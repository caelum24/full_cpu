module array_divider_32b(Q, data_operandA, data_operandB);

    input [31:0] data_operandA, data_operandB;
    // input clock, ctrl_DIV;
    output [31:0] Q;
    // output data_resultRDY;

    wire [62:0] dividend;
    wire [31:0] divisor;
    wire [31:0] div_result;

    //TODO: add registers to store the input values
    //TODO: add clock delay and clock+ctrl_DIV to put together the dataRDY value properly
    //TODO: make dataRDY instant if we have an exception
    
    // assign divisor = data_operandB;
    // assign dividend[31:0] = data_operandA; //replace with output of negating maybe
    
    //negating data_operandA
    wire [31:0] not_A;
    wire isNotEqual_A, isLessThan_A, sub_overflow_A;
    sub_32bit negatorA(not_A, isNotEqual_A, isLessThan_A, sub_overflow_A, 32'b0, data_operandA);
    assign dividend[31:0] = data_operandA[31] ? not_A : data_operandA;
    assign dividend[62:32] = 31'b0;

    //negating data_operandB
    wire [31:0] not_B;
    wire isNotEqual_B, isLessThan_B, sub_overflow_B;
    sub_32bit negatorB(not_B, isNotEqual_B, isLessThan_B, sub_overflow_B, 32'b0, data_operandB);
    assign divisor = data_operandB[31] ? not_B : data_operandB;

    //negating at the end
    wire negator;
    xor (negator, data_operandA[31], data_operandB[31]);
    wire [31:0] not_result;
    wire isNotEqual_o, isLessThan_o, sub_overflow_o;
    sub_32bit negatorC(not_result, isNotEqual_o, isLessThan_o, sub_overflow_o, 32'b0, div_result);
    assign Q = negator ? not_result : div_result;


    wire c_0_0, c_0_1, c_0_2, c_0_3, c_0_4, c_0_5, c_0_6, c_0_7, c_0_8, c_0_9, c_0_10, c_0_11, c_0_12, c_0_13, c_0_14, c_0_15, c_0_16, c_0_17, c_0_18, c_0_19, c_0_20, c_0_21, c_0_22, c_0_23, c_0_24, c_0_25, c_0_26, c_0_27, c_0_28, c_0_29, c_0_30, c_0_31;
    wire empty0, s_0_1, s_0_2, s_0_3, s_0_4, s_0_5, s_0_6, s_0_7, s_0_8, s_0_9, s_0_10, s_0_11, s_0_12, s_0_13, s_0_14, s_0_15, s_0_16, s_0_17, s_0_18, s_0_19, s_0_20, s_0_21, s_0_22, s_0_23, s_0_24, s_0_25, s_0_26, s_0_27, s_0_28, s_0_29, s_0_30, s_0_31;
    divider_cell cell_0_0(empty0, c_0_0, divisor[31], dividend[62], c_0_1, 1'b1);
    divider_cell cell_0_1(s_0_1, c_0_1, divisor[30], dividend[61], c_0_2, 1'b1);
    divider_cell cell_0_2(s_0_2, c_0_2, divisor[29], dividend[60], c_0_3, 1'b1);
    divider_cell cell_0_3(s_0_3, c_0_3, divisor[28], dividend[59], c_0_4, 1'b1);
    divider_cell cell_0_4(s_0_4, c_0_4, divisor[27], dividend[58], c_0_5, 1'b1);
    divider_cell cell_0_5(s_0_5, c_0_5, divisor[26], dividend[57], c_0_6, 1'b1);
    divider_cell cell_0_6(s_0_6, c_0_6, divisor[25], dividend[56], c_0_7, 1'b1);
    divider_cell cell_0_7(s_0_7, c_0_7, divisor[24], dividend[55], c_0_8, 1'b1);
    divider_cell cell_0_8(s_0_8, c_0_8, divisor[23], dividend[54], c_0_9, 1'b1);
    divider_cell cell_0_9(s_0_9, c_0_9, divisor[22], dividend[53], c_0_10, 1'b1);
    divider_cell cell_0_10(s_0_10, c_0_10, divisor[21], dividend[52], c_0_11, 1'b1);
    divider_cell cell_0_11(s_0_11, c_0_11, divisor[20], dividend[51], c_0_12, 1'b1);
    divider_cell cell_0_12(s_0_12, c_0_12, divisor[19], dividend[50], c_0_13, 1'b1);
    divider_cell cell_0_13(s_0_13, c_0_13, divisor[18], dividend[49], c_0_14, 1'b1);
    divider_cell cell_0_14(s_0_14, c_0_14, divisor[17], dividend[48], c_0_15, 1'b1);
    divider_cell cell_0_15(s_0_15, c_0_15, divisor[16], dividend[47], c_0_16, 1'b1);
    divider_cell cell_0_16(s_0_16, c_0_16, divisor[15], dividend[46], c_0_17, 1'b1);
    divider_cell cell_0_17(s_0_17, c_0_17, divisor[14], dividend[45], c_0_18, 1'b1);
    divider_cell cell_0_18(s_0_18, c_0_18, divisor[13], dividend[44], c_0_19, 1'b1);
    divider_cell cell_0_19(s_0_19, c_0_19, divisor[12], dividend[43], c_0_20, 1'b1);
    divider_cell cell_0_20(s_0_20, c_0_20, divisor[11], dividend[42], c_0_21, 1'b1);
    divider_cell cell_0_21(s_0_21, c_0_21, divisor[10], dividend[41], c_0_22, 1'b1);
    divider_cell cell_0_22(s_0_22, c_0_22, divisor[9], dividend[40], c_0_23, 1'b1);
    divider_cell cell_0_23(s_0_23, c_0_23, divisor[8], dividend[39], c_0_24, 1'b1);
    divider_cell cell_0_24(s_0_24, c_0_24, divisor[7], dividend[38], c_0_25, 1'b1);
    divider_cell cell_0_25(s_0_25, c_0_25, divisor[6], dividend[37], c_0_26, 1'b1);
    divider_cell cell_0_26(s_0_26, c_0_26, divisor[5], dividend[36], c_0_27, 1'b1);
    divider_cell cell_0_27(s_0_27, c_0_27, divisor[4], dividend[35], c_0_28, 1'b1);
    divider_cell cell_0_28(s_0_28, c_0_28, divisor[3], dividend[34], c_0_29, 1'b1);
    divider_cell cell_0_29(s_0_29, c_0_29, divisor[2], dividend[33], c_0_30, 1'b1);
    divider_cell cell_0_30(s_0_30, c_0_30, divisor[1], dividend[32], c_0_31, 1'b1);
    divider_cell cell_0_31(s_0_31, c_0_31, divisor[0], dividend[31], 1'b1, 1'b1);
    assign div_result[31] = c_0_0;
    wire c_1_1, c_1_2, c_1_3, c_1_4, c_1_5, c_1_6, c_1_7, c_1_8, c_1_9, c_1_10, c_1_11, c_1_12, c_1_13, c_1_14, c_1_15, c_1_16, c_1_17, c_1_18, c_1_19, c_1_20, c_1_21, c_1_22, c_1_23, c_1_24, c_1_25, c_1_26, c_1_27, c_1_28, c_1_29, c_1_30, c_1_31, c_1_32;
    wire empty1, s_1_2, s_1_3, s_1_4, s_1_5, s_1_6, s_1_7, s_1_8, s_1_9, s_1_10, s_1_11, s_1_12, s_1_13, s_1_14, s_1_15, s_1_16, s_1_17, s_1_18, s_1_19, s_1_20, s_1_21, s_1_22, s_1_23, s_1_24, s_1_25, s_1_26, s_1_27, s_1_28, s_1_29, s_1_30, s_1_31, s_1_32;
    divider_cell cell_1_1(empty1, c_1_1, divisor[31], s_0_1, c_1_2, c_0_0);
    divider_cell cell_1_2(s_1_2, c_1_2, divisor[30], s_0_2, c_1_3, c_0_0);
    divider_cell cell_1_3(s_1_3, c_1_3, divisor[29], s_0_3, c_1_4, c_0_0);
    divider_cell cell_1_4(s_1_4, c_1_4, divisor[28], s_0_4, c_1_5, c_0_0);
    divider_cell cell_1_5(s_1_5, c_1_5, divisor[27], s_0_5, c_1_6, c_0_0);
    divider_cell cell_1_6(s_1_6, c_1_6, divisor[26], s_0_6, c_1_7, c_0_0);
    divider_cell cell_1_7(s_1_7, c_1_7, divisor[25], s_0_7, c_1_8, c_0_0);
    divider_cell cell_1_8(s_1_8, c_1_8, divisor[24], s_0_8, c_1_9, c_0_0);
    divider_cell cell_1_9(s_1_9, c_1_9, divisor[23], s_0_9, c_1_10, c_0_0);
    divider_cell cell_1_10(s_1_10, c_1_10, divisor[22], s_0_10, c_1_11, c_0_0);
    divider_cell cell_1_11(s_1_11, c_1_11, divisor[21], s_0_11, c_1_12, c_0_0);
    divider_cell cell_1_12(s_1_12, c_1_12, divisor[20], s_0_12, c_1_13, c_0_0);
    divider_cell cell_1_13(s_1_13, c_1_13, divisor[19], s_0_13, c_1_14, c_0_0);
    divider_cell cell_1_14(s_1_14, c_1_14, divisor[18], s_0_14, c_1_15, c_0_0);
    divider_cell cell_1_15(s_1_15, c_1_15, divisor[17], s_0_15, c_1_16, c_0_0);
    divider_cell cell_1_16(s_1_16, c_1_16, divisor[16], s_0_16, c_1_17, c_0_0);
    divider_cell cell_1_17(s_1_17, c_1_17, divisor[15], s_0_17, c_1_18, c_0_0);
    divider_cell cell_1_18(s_1_18, c_1_18, divisor[14], s_0_18, c_1_19, c_0_0);
    divider_cell cell_1_19(s_1_19, c_1_19, divisor[13], s_0_19, c_1_20, c_0_0);
    divider_cell cell_1_20(s_1_20, c_1_20, divisor[12], s_0_20, c_1_21, c_0_0);
    divider_cell cell_1_21(s_1_21, c_1_21, divisor[11], s_0_21, c_1_22, c_0_0);
    divider_cell cell_1_22(s_1_22, c_1_22, divisor[10], s_0_22, c_1_23, c_0_0);
    divider_cell cell_1_23(s_1_23, c_1_23, divisor[9], s_0_23, c_1_24, c_0_0);
    divider_cell cell_1_24(s_1_24, c_1_24, divisor[8], s_0_24, c_1_25, c_0_0);
    divider_cell cell_1_25(s_1_25, c_1_25, divisor[7], s_0_25, c_1_26, c_0_0);
    divider_cell cell_1_26(s_1_26, c_1_26, divisor[6], s_0_26, c_1_27, c_0_0);
    divider_cell cell_1_27(s_1_27, c_1_27, divisor[5], s_0_27, c_1_28, c_0_0);
    divider_cell cell_1_28(s_1_28, c_1_28, divisor[4], s_0_28, c_1_29, c_0_0);
    divider_cell cell_1_29(s_1_29, c_1_29, divisor[3], s_0_29, c_1_30, c_0_0);
    divider_cell cell_1_30(s_1_30, c_1_30, divisor[2], s_0_30, c_1_31, c_0_0);
    divider_cell cell_1_31(s_1_31, c_1_31, divisor[1], s_0_31, c_1_32, c_0_0);
    divider_cell cell_1_32(s_1_32, c_1_32, divisor[0], dividend[30], c_0_0, c_0_0);
    assign div_result[30] = c_1_1;
    wire c_2_2, c_2_3, c_2_4, c_2_5, c_2_6, c_2_7, c_2_8, c_2_9, c_2_10, c_2_11, c_2_12, c_2_13, c_2_14, c_2_15, c_2_16, c_2_17, c_2_18, c_2_19, c_2_20, c_2_21, c_2_22, c_2_23, c_2_24, c_2_25, c_2_26, c_2_27, c_2_28, c_2_29, c_2_30, c_2_31, c_2_32, c_2_33;
    wire empty2, s_2_3, s_2_4, s_2_5, s_2_6, s_2_7, s_2_8, s_2_9, s_2_10, s_2_11, s_2_12, s_2_13, s_2_14, s_2_15, s_2_16, s_2_17, s_2_18, s_2_19, s_2_20, s_2_21, s_2_22, s_2_23, s_2_24, s_2_25, s_2_26, s_2_27, s_2_28, s_2_29, s_2_30, s_2_31, s_2_32, s_2_33;
    divider_cell cell_2_2(empty2, c_2_2, divisor[31], s_1_2, c_2_3, c_1_1);
    divider_cell cell_2_3(s_2_3, c_2_3, divisor[30], s_1_3, c_2_4, c_1_1);
    divider_cell cell_2_4(s_2_4, c_2_4, divisor[29], s_1_4, c_2_5, c_1_1);
    divider_cell cell_2_5(s_2_5, c_2_5, divisor[28], s_1_5, c_2_6, c_1_1);
    divider_cell cell_2_6(s_2_6, c_2_6, divisor[27], s_1_6, c_2_7, c_1_1);
    divider_cell cell_2_7(s_2_7, c_2_7, divisor[26], s_1_7, c_2_8, c_1_1);
    divider_cell cell_2_8(s_2_8, c_2_8, divisor[25], s_1_8, c_2_9, c_1_1);
    divider_cell cell_2_9(s_2_9, c_2_9, divisor[24], s_1_9, c_2_10, c_1_1);
    divider_cell cell_2_10(s_2_10, c_2_10, divisor[23], s_1_10, c_2_11, c_1_1);
    divider_cell cell_2_11(s_2_11, c_2_11, divisor[22], s_1_11, c_2_12, c_1_1);
    divider_cell cell_2_12(s_2_12, c_2_12, divisor[21], s_1_12, c_2_13, c_1_1);
    divider_cell cell_2_13(s_2_13, c_2_13, divisor[20], s_1_13, c_2_14, c_1_1);
    divider_cell cell_2_14(s_2_14, c_2_14, divisor[19], s_1_14, c_2_15, c_1_1);
    divider_cell cell_2_15(s_2_15, c_2_15, divisor[18], s_1_15, c_2_16, c_1_1);
    divider_cell cell_2_16(s_2_16, c_2_16, divisor[17], s_1_16, c_2_17, c_1_1);
    divider_cell cell_2_17(s_2_17, c_2_17, divisor[16], s_1_17, c_2_18, c_1_1);
    divider_cell cell_2_18(s_2_18, c_2_18, divisor[15], s_1_18, c_2_19, c_1_1);
    divider_cell cell_2_19(s_2_19, c_2_19, divisor[14], s_1_19, c_2_20, c_1_1);
    divider_cell cell_2_20(s_2_20, c_2_20, divisor[13], s_1_20, c_2_21, c_1_1);
    divider_cell cell_2_21(s_2_21, c_2_21, divisor[12], s_1_21, c_2_22, c_1_1);
    divider_cell cell_2_22(s_2_22, c_2_22, divisor[11], s_1_22, c_2_23, c_1_1);
    divider_cell cell_2_23(s_2_23, c_2_23, divisor[10], s_1_23, c_2_24, c_1_1);
    divider_cell cell_2_24(s_2_24, c_2_24, divisor[9], s_1_24, c_2_25, c_1_1);
    divider_cell cell_2_25(s_2_25, c_2_25, divisor[8], s_1_25, c_2_26, c_1_1);
    divider_cell cell_2_26(s_2_26, c_2_26, divisor[7], s_1_26, c_2_27, c_1_1);
    divider_cell cell_2_27(s_2_27, c_2_27, divisor[6], s_1_27, c_2_28, c_1_1);
    divider_cell cell_2_28(s_2_28, c_2_28, divisor[5], s_1_28, c_2_29, c_1_1);
    divider_cell cell_2_29(s_2_29, c_2_29, divisor[4], s_1_29, c_2_30, c_1_1);
    divider_cell cell_2_30(s_2_30, c_2_30, divisor[3], s_1_30, c_2_31, c_1_1);
    divider_cell cell_2_31(s_2_31, c_2_31, divisor[2], s_1_31, c_2_32, c_1_1);
    divider_cell cell_2_32(s_2_32, c_2_32, divisor[1], s_1_32, c_2_33, c_1_1);
    divider_cell cell_2_33(s_2_33, c_2_33, divisor[0], dividend[29], c_1_1, c_1_1);
    assign div_result[29] = c_2_2;
    wire c_3_3, c_3_4, c_3_5, c_3_6, c_3_7, c_3_8, c_3_9, c_3_10, c_3_11, c_3_12, c_3_13, c_3_14, c_3_15, c_3_16, c_3_17, c_3_18, c_3_19, c_3_20, c_3_21, c_3_22, c_3_23, c_3_24, c_3_25, c_3_26, c_3_27, c_3_28, c_3_29, c_3_30, c_3_31, c_3_32, c_3_33, c_3_34;
    wire empty3, s_3_4, s_3_5, s_3_6, s_3_7, s_3_8, s_3_9, s_3_10, s_3_11, s_3_12, s_3_13, s_3_14, s_3_15, s_3_16, s_3_17, s_3_18, s_3_19, s_3_20, s_3_21, s_3_22, s_3_23, s_3_24, s_3_25, s_3_26, s_3_27, s_3_28, s_3_29, s_3_30, s_3_31, s_3_32, s_3_33, s_3_34;
    divider_cell cell_3_3(empty3, c_3_3, divisor[31], s_2_3, c_3_4, c_2_2);
    divider_cell cell_3_4(s_3_4, c_3_4, divisor[30], s_2_4, c_3_5, c_2_2);
    divider_cell cell_3_5(s_3_5, c_3_5, divisor[29], s_2_5, c_3_6, c_2_2);
    divider_cell cell_3_6(s_3_6, c_3_6, divisor[28], s_2_6, c_3_7, c_2_2);
    divider_cell cell_3_7(s_3_7, c_3_7, divisor[27], s_2_7, c_3_8, c_2_2);
    divider_cell cell_3_8(s_3_8, c_3_8, divisor[26], s_2_8, c_3_9, c_2_2);
    divider_cell cell_3_9(s_3_9, c_3_9, divisor[25], s_2_9, c_3_10, c_2_2);
    divider_cell cell_3_10(s_3_10, c_3_10, divisor[24], s_2_10, c_3_11, c_2_2);
    divider_cell cell_3_11(s_3_11, c_3_11, divisor[23], s_2_11, c_3_12, c_2_2);
    divider_cell cell_3_12(s_3_12, c_3_12, divisor[22], s_2_12, c_3_13, c_2_2);
    divider_cell cell_3_13(s_3_13, c_3_13, divisor[21], s_2_13, c_3_14, c_2_2);
    divider_cell cell_3_14(s_3_14, c_3_14, divisor[20], s_2_14, c_3_15, c_2_2);
    divider_cell cell_3_15(s_3_15, c_3_15, divisor[19], s_2_15, c_3_16, c_2_2);
    divider_cell cell_3_16(s_3_16, c_3_16, divisor[18], s_2_16, c_3_17, c_2_2);
    divider_cell cell_3_17(s_3_17, c_3_17, divisor[17], s_2_17, c_3_18, c_2_2);
    divider_cell cell_3_18(s_3_18, c_3_18, divisor[16], s_2_18, c_3_19, c_2_2);
    divider_cell cell_3_19(s_3_19, c_3_19, divisor[15], s_2_19, c_3_20, c_2_2);
    divider_cell cell_3_20(s_3_20, c_3_20, divisor[14], s_2_20, c_3_21, c_2_2);
    divider_cell cell_3_21(s_3_21, c_3_21, divisor[13], s_2_21, c_3_22, c_2_2);
    divider_cell cell_3_22(s_3_22, c_3_22, divisor[12], s_2_22, c_3_23, c_2_2);
    divider_cell cell_3_23(s_3_23, c_3_23, divisor[11], s_2_23, c_3_24, c_2_2);
    divider_cell cell_3_24(s_3_24, c_3_24, divisor[10], s_2_24, c_3_25, c_2_2);
    divider_cell cell_3_25(s_3_25, c_3_25, divisor[9], s_2_25, c_3_26, c_2_2);
    divider_cell cell_3_26(s_3_26, c_3_26, divisor[8], s_2_26, c_3_27, c_2_2);
    divider_cell cell_3_27(s_3_27, c_3_27, divisor[7], s_2_27, c_3_28, c_2_2);
    divider_cell cell_3_28(s_3_28, c_3_28, divisor[6], s_2_28, c_3_29, c_2_2);
    divider_cell cell_3_29(s_3_29, c_3_29, divisor[5], s_2_29, c_3_30, c_2_2);
    divider_cell cell_3_30(s_3_30, c_3_30, divisor[4], s_2_30, c_3_31, c_2_2);
    divider_cell cell_3_31(s_3_31, c_3_31, divisor[3], s_2_31, c_3_32, c_2_2);
    divider_cell cell_3_32(s_3_32, c_3_32, divisor[2], s_2_32, c_3_33, c_2_2);
    divider_cell cell_3_33(s_3_33, c_3_33, divisor[1], s_2_33, c_3_34, c_2_2);
    divider_cell cell_3_34(s_3_34, c_3_34, divisor[0], dividend[28], c_2_2, c_2_2);
    assign div_result[28] = c_3_3;
    wire c_4_4, c_4_5, c_4_6, c_4_7, c_4_8, c_4_9, c_4_10, c_4_11, c_4_12, c_4_13, c_4_14, c_4_15, c_4_16, c_4_17, c_4_18, c_4_19, c_4_20, c_4_21, c_4_22, c_4_23, c_4_24, c_4_25, c_4_26, c_4_27, c_4_28, c_4_29, c_4_30, c_4_31, c_4_32, c_4_33, c_4_34, c_4_35;
    wire empty4, s_4_5, s_4_6, s_4_7, s_4_8, s_4_9, s_4_10, s_4_11, s_4_12, s_4_13, s_4_14, s_4_15, s_4_16, s_4_17, s_4_18, s_4_19, s_4_20, s_4_21, s_4_22, s_4_23, s_4_24, s_4_25, s_4_26, s_4_27, s_4_28, s_4_29, s_4_30, s_4_31, s_4_32, s_4_33, s_4_34, s_4_35;
    divider_cell cell_4_4(empty4, c_4_4, divisor[31], s_3_4, c_4_5, c_3_3);
    divider_cell cell_4_5(s_4_5, c_4_5, divisor[30], s_3_5, c_4_6, c_3_3);
    divider_cell cell_4_6(s_4_6, c_4_6, divisor[29], s_3_6, c_4_7, c_3_3);
    divider_cell cell_4_7(s_4_7, c_4_7, divisor[28], s_3_7, c_4_8, c_3_3);
    divider_cell cell_4_8(s_4_8, c_4_8, divisor[27], s_3_8, c_4_9, c_3_3);
    divider_cell cell_4_9(s_4_9, c_4_9, divisor[26], s_3_9, c_4_10, c_3_3);
    divider_cell cell_4_10(s_4_10, c_4_10, divisor[25], s_3_10, c_4_11, c_3_3);
    divider_cell cell_4_11(s_4_11, c_4_11, divisor[24], s_3_11, c_4_12, c_3_3);
    divider_cell cell_4_12(s_4_12, c_4_12, divisor[23], s_3_12, c_4_13, c_3_3);
    divider_cell cell_4_13(s_4_13, c_4_13, divisor[22], s_3_13, c_4_14, c_3_3);
    divider_cell cell_4_14(s_4_14, c_4_14, divisor[21], s_3_14, c_4_15, c_3_3);
    divider_cell cell_4_15(s_4_15, c_4_15, divisor[20], s_3_15, c_4_16, c_3_3);
    divider_cell cell_4_16(s_4_16, c_4_16, divisor[19], s_3_16, c_4_17, c_3_3);
    divider_cell cell_4_17(s_4_17, c_4_17, divisor[18], s_3_17, c_4_18, c_3_3);
    divider_cell cell_4_18(s_4_18, c_4_18, divisor[17], s_3_18, c_4_19, c_3_3);
    divider_cell cell_4_19(s_4_19, c_4_19, divisor[16], s_3_19, c_4_20, c_3_3);
    divider_cell cell_4_20(s_4_20, c_4_20, divisor[15], s_3_20, c_4_21, c_3_3);
    divider_cell cell_4_21(s_4_21, c_4_21, divisor[14], s_3_21, c_4_22, c_3_3);
    divider_cell cell_4_22(s_4_22, c_4_22, divisor[13], s_3_22, c_4_23, c_3_3);
    divider_cell cell_4_23(s_4_23, c_4_23, divisor[12], s_3_23, c_4_24, c_3_3);
    divider_cell cell_4_24(s_4_24, c_4_24, divisor[11], s_3_24, c_4_25, c_3_3);
    divider_cell cell_4_25(s_4_25, c_4_25, divisor[10], s_3_25, c_4_26, c_3_3);
    divider_cell cell_4_26(s_4_26, c_4_26, divisor[9], s_3_26, c_4_27, c_3_3);
    divider_cell cell_4_27(s_4_27, c_4_27, divisor[8], s_3_27, c_4_28, c_3_3);
    divider_cell cell_4_28(s_4_28, c_4_28, divisor[7], s_3_28, c_4_29, c_3_3);
    divider_cell cell_4_29(s_4_29, c_4_29, divisor[6], s_3_29, c_4_30, c_3_3);
    divider_cell cell_4_30(s_4_30, c_4_30, divisor[5], s_3_30, c_4_31, c_3_3);
    divider_cell cell_4_31(s_4_31, c_4_31, divisor[4], s_3_31, c_4_32, c_3_3);
    divider_cell cell_4_32(s_4_32, c_4_32, divisor[3], s_3_32, c_4_33, c_3_3);
    divider_cell cell_4_33(s_4_33, c_4_33, divisor[2], s_3_33, c_4_34, c_3_3);
    divider_cell cell_4_34(s_4_34, c_4_34, divisor[1], s_3_34, c_4_35, c_3_3);
    divider_cell cell_4_35(s_4_35, c_4_35, divisor[0], dividend[27], c_3_3, c_3_3);
    assign div_result[27] = c_4_4;
    wire c_5_5, c_5_6, c_5_7, c_5_8, c_5_9, c_5_10, c_5_11, c_5_12, c_5_13, c_5_14, c_5_15, c_5_16, c_5_17, c_5_18, c_5_19, c_5_20, c_5_21, c_5_22, c_5_23, c_5_24, c_5_25, c_5_26, c_5_27, c_5_28, c_5_29, c_5_30, c_5_31, c_5_32, c_5_33, c_5_34, c_5_35, c_5_36;
    wire empty5, s_5_6, s_5_7, s_5_8, s_5_9, s_5_10, s_5_11, s_5_12, s_5_13, s_5_14, s_5_15, s_5_16, s_5_17, s_5_18, s_5_19, s_5_20, s_5_21, s_5_22, s_5_23, s_5_24, s_5_25, s_5_26, s_5_27, s_5_28, s_5_29, s_5_30, s_5_31, s_5_32, s_5_33, s_5_34, s_5_35, s_5_36;
    divider_cell cell_5_5(empty5, c_5_5, divisor[31], s_4_5, c_5_6, c_4_4);
    divider_cell cell_5_6(s_5_6, c_5_6, divisor[30], s_4_6, c_5_7, c_4_4);
    divider_cell cell_5_7(s_5_7, c_5_7, divisor[29], s_4_7, c_5_8, c_4_4);
    divider_cell cell_5_8(s_5_8, c_5_8, divisor[28], s_4_8, c_5_9, c_4_4);
    divider_cell cell_5_9(s_5_9, c_5_9, divisor[27], s_4_9, c_5_10, c_4_4);
    divider_cell cell_5_10(s_5_10, c_5_10, divisor[26], s_4_10, c_5_11, c_4_4);
    divider_cell cell_5_11(s_5_11, c_5_11, divisor[25], s_4_11, c_5_12, c_4_4);
    divider_cell cell_5_12(s_5_12, c_5_12, divisor[24], s_4_12, c_5_13, c_4_4);
    divider_cell cell_5_13(s_5_13, c_5_13, divisor[23], s_4_13, c_5_14, c_4_4);
    divider_cell cell_5_14(s_5_14, c_5_14, divisor[22], s_4_14, c_5_15, c_4_4);
    divider_cell cell_5_15(s_5_15, c_5_15, divisor[21], s_4_15, c_5_16, c_4_4);
    divider_cell cell_5_16(s_5_16, c_5_16, divisor[20], s_4_16, c_5_17, c_4_4);
    divider_cell cell_5_17(s_5_17, c_5_17, divisor[19], s_4_17, c_5_18, c_4_4);
    divider_cell cell_5_18(s_5_18, c_5_18, divisor[18], s_4_18, c_5_19, c_4_4);
    divider_cell cell_5_19(s_5_19, c_5_19, divisor[17], s_4_19, c_5_20, c_4_4);
    divider_cell cell_5_20(s_5_20, c_5_20, divisor[16], s_4_20, c_5_21, c_4_4);
    divider_cell cell_5_21(s_5_21, c_5_21, divisor[15], s_4_21, c_5_22, c_4_4);
    divider_cell cell_5_22(s_5_22, c_5_22, divisor[14], s_4_22, c_5_23, c_4_4);
    divider_cell cell_5_23(s_5_23, c_5_23, divisor[13], s_4_23, c_5_24, c_4_4);
    divider_cell cell_5_24(s_5_24, c_5_24, divisor[12], s_4_24, c_5_25, c_4_4);
    divider_cell cell_5_25(s_5_25, c_5_25, divisor[11], s_4_25, c_5_26, c_4_4);
    divider_cell cell_5_26(s_5_26, c_5_26, divisor[10], s_4_26, c_5_27, c_4_4);
    divider_cell cell_5_27(s_5_27, c_5_27, divisor[9], s_4_27, c_5_28, c_4_4);
    divider_cell cell_5_28(s_5_28, c_5_28, divisor[8], s_4_28, c_5_29, c_4_4);
    divider_cell cell_5_29(s_5_29, c_5_29, divisor[7], s_4_29, c_5_30, c_4_4);
    divider_cell cell_5_30(s_5_30, c_5_30, divisor[6], s_4_30, c_5_31, c_4_4);
    divider_cell cell_5_31(s_5_31, c_5_31, divisor[5], s_4_31, c_5_32, c_4_4);
    divider_cell cell_5_32(s_5_32, c_5_32, divisor[4], s_4_32, c_5_33, c_4_4);
    divider_cell cell_5_33(s_5_33, c_5_33, divisor[3], s_4_33, c_5_34, c_4_4);
    divider_cell cell_5_34(s_5_34, c_5_34, divisor[2], s_4_34, c_5_35, c_4_4);
    divider_cell cell_5_35(s_5_35, c_5_35, divisor[1], s_4_35, c_5_36, c_4_4);
    divider_cell cell_5_36(s_5_36, c_5_36, divisor[0], dividend[26], c_4_4, c_4_4);
    assign div_result[26] = c_5_5;
    wire c_6_6, c_6_7, c_6_8, c_6_9, c_6_10, c_6_11, c_6_12, c_6_13, c_6_14, c_6_15, c_6_16, c_6_17, c_6_18, c_6_19, c_6_20, c_6_21, c_6_22, c_6_23, c_6_24, c_6_25, c_6_26, c_6_27, c_6_28, c_6_29, c_6_30, c_6_31, c_6_32, c_6_33, c_6_34, c_6_35, c_6_36, c_6_37;
    wire empty6, s_6_7, s_6_8, s_6_9, s_6_10, s_6_11, s_6_12, s_6_13, s_6_14, s_6_15, s_6_16, s_6_17, s_6_18, s_6_19, s_6_20, s_6_21, s_6_22, s_6_23, s_6_24, s_6_25, s_6_26, s_6_27, s_6_28, s_6_29, s_6_30, s_6_31, s_6_32, s_6_33, s_6_34, s_6_35, s_6_36, s_6_37;
    divider_cell cell_6_6(empty6, c_6_6, divisor[31], s_5_6, c_6_7, c_5_5);
    divider_cell cell_6_7(s_6_7, c_6_7, divisor[30], s_5_7, c_6_8, c_5_5);
    divider_cell cell_6_8(s_6_8, c_6_8, divisor[29], s_5_8, c_6_9, c_5_5);
    divider_cell cell_6_9(s_6_9, c_6_9, divisor[28], s_5_9, c_6_10, c_5_5);
    divider_cell cell_6_10(s_6_10, c_6_10, divisor[27], s_5_10, c_6_11, c_5_5);
    divider_cell cell_6_11(s_6_11, c_6_11, divisor[26], s_5_11, c_6_12, c_5_5);
    divider_cell cell_6_12(s_6_12, c_6_12, divisor[25], s_5_12, c_6_13, c_5_5);
    divider_cell cell_6_13(s_6_13, c_6_13, divisor[24], s_5_13, c_6_14, c_5_5);
    divider_cell cell_6_14(s_6_14, c_6_14, divisor[23], s_5_14, c_6_15, c_5_5);
    divider_cell cell_6_15(s_6_15, c_6_15, divisor[22], s_5_15, c_6_16, c_5_5);
    divider_cell cell_6_16(s_6_16, c_6_16, divisor[21], s_5_16, c_6_17, c_5_5);
    divider_cell cell_6_17(s_6_17, c_6_17, divisor[20], s_5_17, c_6_18, c_5_5);
    divider_cell cell_6_18(s_6_18, c_6_18, divisor[19], s_5_18, c_6_19, c_5_5);
    divider_cell cell_6_19(s_6_19, c_6_19, divisor[18], s_5_19, c_6_20, c_5_5);
    divider_cell cell_6_20(s_6_20, c_6_20, divisor[17], s_5_20, c_6_21, c_5_5);
    divider_cell cell_6_21(s_6_21, c_6_21, divisor[16], s_5_21, c_6_22, c_5_5);
    divider_cell cell_6_22(s_6_22, c_6_22, divisor[15], s_5_22, c_6_23, c_5_5);
    divider_cell cell_6_23(s_6_23, c_6_23, divisor[14], s_5_23, c_6_24, c_5_5);
    divider_cell cell_6_24(s_6_24, c_6_24, divisor[13], s_5_24, c_6_25, c_5_5);
    divider_cell cell_6_25(s_6_25, c_6_25, divisor[12], s_5_25, c_6_26, c_5_5);
    divider_cell cell_6_26(s_6_26, c_6_26, divisor[11], s_5_26, c_6_27, c_5_5);
    divider_cell cell_6_27(s_6_27, c_6_27, divisor[10], s_5_27, c_6_28, c_5_5);
    divider_cell cell_6_28(s_6_28, c_6_28, divisor[9], s_5_28, c_6_29, c_5_5);
    divider_cell cell_6_29(s_6_29, c_6_29, divisor[8], s_5_29, c_6_30, c_5_5);
    divider_cell cell_6_30(s_6_30, c_6_30, divisor[7], s_5_30, c_6_31, c_5_5);
    divider_cell cell_6_31(s_6_31, c_6_31, divisor[6], s_5_31, c_6_32, c_5_5);
    divider_cell cell_6_32(s_6_32, c_6_32, divisor[5], s_5_32, c_6_33, c_5_5);
    divider_cell cell_6_33(s_6_33, c_6_33, divisor[4], s_5_33, c_6_34, c_5_5);
    divider_cell cell_6_34(s_6_34, c_6_34, divisor[3], s_5_34, c_6_35, c_5_5);
    divider_cell cell_6_35(s_6_35, c_6_35, divisor[2], s_5_35, c_6_36, c_5_5);
    divider_cell cell_6_36(s_6_36, c_6_36, divisor[1], s_5_36, c_6_37, c_5_5);
    divider_cell cell_6_37(s_6_37, c_6_37, divisor[0], dividend[25], c_5_5, c_5_5);
    assign div_result[25] = c_6_6;
    wire c_7_7, c_7_8, c_7_9, c_7_10, c_7_11, c_7_12, c_7_13, c_7_14, c_7_15, c_7_16, c_7_17, c_7_18, c_7_19, c_7_20, c_7_21, c_7_22, c_7_23, c_7_24, c_7_25, c_7_26, c_7_27, c_7_28, c_7_29, c_7_30, c_7_31, c_7_32, c_7_33, c_7_34, c_7_35, c_7_36, c_7_37, c_7_38;
    wire empty7, s_7_8, s_7_9, s_7_10, s_7_11, s_7_12, s_7_13, s_7_14, s_7_15, s_7_16, s_7_17, s_7_18, s_7_19, s_7_20, s_7_21, s_7_22, s_7_23, s_7_24, s_7_25, s_7_26, s_7_27, s_7_28, s_7_29, s_7_30, s_7_31, s_7_32, s_7_33, s_7_34, s_7_35, s_7_36, s_7_37, s_7_38;
    divider_cell cell_7_7(empty7, c_7_7, divisor[31], s_6_7, c_7_8, c_6_6);
    divider_cell cell_7_8(s_7_8, c_7_8, divisor[30], s_6_8, c_7_9, c_6_6);
    divider_cell cell_7_9(s_7_9, c_7_9, divisor[29], s_6_9, c_7_10, c_6_6);
    divider_cell cell_7_10(s_7_10, c_7_10, divisor[28], s_6_10, c_7_11, c_6_6);
    divider_cell cell_7_11(s_7_11, c_7_11, divisor[27], s_6_11, c_7_12, c_6_6);
    divider_cell cell_7_12(s_7_12, c_7_12, divisor[26], s_6_12, c_7_13, c_6_6);
    divider_cell cell_7_13(s_7_13, c_7_13, divisor[25], s_6_13, c_7_14, c_6_6);
    divider_cell cell_7_14(s_7_14, c_7_14, divisor[24], s_6_14, c_7_15, c_6_6);
    divider_cell cell_7_15(s_7_15, c_7_15, divisor[23], s_6_15, c_7_16, c_6_6);
    divider_cell cell_7_16(s_7_16, c_7_16, divisor[22], s_6_16, c_7_17, c_6_6);
    divider_cell cell_7_17(s_7_17, c_7_17, divisor[21], s_6_17, c_7_18, c_6_6);
    divider_cell cell_7_18(s_7_18, c_7_18, divisor[20], s_6_18, c_7_19, c_6_6);
    divider_cell cell_7_19(s_7_19, c_7_19, divisor[19], s_6_19, c_7_20, c_6_6);
    divider_cell cell_7_20(s_7_20, c_7_20, divisor[18], s_6_20, c_7_21, c_6_6);
    divider_cell cell_7_21(s_7_21, c_7_21, divisor[17], s_6_21, c_7_22, c_6_6);
    divider_cell cell_7_22(s_7_22, c_7_22, divisor[16], s_6_22, c_7_23, c_6_6);
    divider_cell cell_7_23(s_7_23, c_7_23, divisor[15], s_6_23, c_7_24, c_6_6);
    divider_cell cell_7_24(s_7_24, c_7_24, divisor[14], s_6_24, c_7_25, c_6_6);
    divider_cell cell_7_25(s_7_25, c_7_25, divisor[13], s_6_25, c_7_26, c_6_6);
    divider_cell cell_7_26(s_7_26, c_7_26, divisor[12], s_6_26, c_7_27, c_6_6);
    divider_cell cell_7_27(s_7_27, c_7_27, divisor[11], s_6_27, c_7_28, c_6_6);
    divider_cell cell_7_28(s_7_28, c_7_28, divisor[10], s_6_28, c_7_29, c_6_6);
    divider_cell cell_7_29(s_7_29, c_7_29, divisor[9], s_6_29, c_7_30, c_6_6);
    divider_cell cell_7_30(s_7_30, c_7_30, divisor[8], s_6_30, c_7_31, c_6_6);
    divider_cell cell_7_31(s_7_31, c_7_31, divisor[7], s_6_31, c_7_32, c_6_6);
    divider_cell cell_7_32(s_7_32, c_7_32, divisor[6], s_6_32, c_7_33, c_6_6);
    divider_cell cell_7_33(s_7_33, c_7_33, divisor[5], s_6_33, c_7_34, c_6_6);
    divider_cell cell_7_34(s_7_34, c_7_34, divisor[4], s_6_34, c_7_35, c_6_6);
    divider_cell cell_7_35(s_7_35, c_7_35, divisor[3], s_6_35, c_7_36, c_6_6);
    divider_cell cell_7_36(s_7_36, c_7_36, divisor[2], s_6_36, c_7_37, c_6_6);
    divider_cell cell_7_37(s_7_37, c_7_37, divisor[1], s_6_37, c_7_38, c_6_6);
    divider_cell cell_7_38(s_7_38, c_7_38, divisor[0], dividend[24], c_6_6, c_6_6);
    assign div_result[24] = c_7_7;
    wire c_8_8, c_8_9, c_8_10, c_8_11, c_8_12, c_8_13, c_8_14, c_8_15, c_8_16, c_8_17, c_8_18, c_8_19, c_8_20, c_8_21, c_8_22, c_8_23, c_8_24, c_8_25, c_8_26, c_8_27, c_8_28, c_8_29, c_8_30, c_8_31, c_8_32, c_8_33, c_8_34, c_8_35, c_8_36, c_8_37, c_8_38, c_8_39;
    wire empty8, s_8_9, s_8_10, s_8_11, s_8_12, s_8_13, s_8_14, s_8_15, s_8_16, s_8_17, s_8_18, s_8_19, s_8_20, s_8_21, s_8_22, s_8_23, s_8_24, s_8_25, s_8_26, s_8_27, s_8_28, s_8_29, s_8_30, s_8_31, s_8_32, s_8_33, s_8_34, s_8_35, s_8_36, s_8_37, s_8_38, s_8_39;
    divider_cell cell_8_8(empty8, c_8_8, divisor[31], s_7_8, c_8_9, c_7_7);
    divider_cell cell_8_9(s_8_9, c_8_9, divisor[30], s_7_9, c_8_10, c_7_7);
    divider_cell cell_8_10(s_8_10, c_8_10, divisor[29], s_7_10, c_8_11, c_7_7);
    divider_cell cell_8_11(s_8_11, c_8_11, divisor[28], s_7_11, c_8_12, c_7_7);
    divider_cell cell_8_12(s_8_12, c_8_12, divisor[27], s_7_12, c_8_13, c_7_7);
    divider_cell cell_8_13(s_8_13, c_8_13, divisor[26], s_7_13, c_8_14, c_7_7);
    divider_cell cell_8_14(s_8_14, c_8_14, divisor[25], s_7_14, c_8_15, c_7_7);
    divider_cell cell_8_15(s_8_15, c_8_15, divisor[24], s_7_15, c_8_16, c_7_7);
    divider_cell cell_8_16(s_8_16, c_8_16, divisor[23], s_7_16, c_8_17, c_7_7);
    divider_cell cell_8_17(s_8_17, c_8_17, divisor[22], s_7_17, c_8_18, c_7_7);
    divider_cell cell_8_18(s_8_18, c_8_18, divisor[21], s_7_18, c_8_19, c_7_7);
    divider_cell cell_8_19(s_8_19, c_8_19, divisor[20], s_7_19, c_8_20, c_7_7);
    divider_cell cell_8_20(s_8_20, c_8_20, divisor[19], s_7_20, c_8_21, c_7_7);
    divider_cell cell_8_21(s_8_21, c_8_21, divisor[18], s_7_21, c_8_22, c_7_7);
    divider_cell cell_8_22(s_8_22, c_8_22, divisor[17], s_7_22, c_8_23, c_7_7);
    divider_cell cell_8_23(s_8_23, c_8_23, divisor[16], s_7_23, c_8_24, c_7_7);
    divider_cell cell_8_24(s_8_24, c_8_24, divisor[15], s_7_24, c_8_25, c_7_7);
    divider_cell cell_8_25(s_8_25, c_8_25, divisor[14], s_7_25, c_8_26, c_7_7);
    divider_cell cell_8_26(s_8_26, c_8_26, divisor[13], s_7_26, c_8_27, c_7_7);
    divider_cell cell_8_27(s_8_27, c_8_27, divisor[12], s_7_27, c_8_28, c_7_7);
    divider_cell cell_8_28(s_8_28, c_8_28, divisor[11], s_7_28, c_8_29, c_7_7);
    divider_cell cell_8_29(s_8_29, c_8_29, divisor[10], s_7_29, c_8_30, c_7_7);
    divider_cell cell_8_30(s_8_30, c_8_30, divisor[9], s_7_30, c_8_31, c_7_7);
    divider_cell cell_8_31(s_8_31, c_8_31, divisor[8], s_7_31, c_8_32, c_7_7);
    divider_cell cell_8_32(s_8_32, c_8_32, divisor[7], s_7_32, c_8_33, c_7_7);
    divider_cell cell_8_33(s_8_33, c_8_33, divisor[6], s_7_33, c_8_34, c_7_7);
    divider_cell cell_8_34(s_8_34, c_8_34, divisor[5], s_7_34, c_8_35, c_7_7);
    divider_cell cell_8_35(s_8_35, c_8_35, divisor[4], s_7_35, c_8_36, c_7_7);
    divider_cell cell_8_36(s_8_36, c_8_36, divisor[3], s_7_36, c_8_37, c_7_7);
    divider_cell cell_8_37(s_8_37, c_8_37, divisor[2], s_7_37, c_8_38, c_7_7);
    divider_cell cell_8_38(s_8_38, c_8_38, divisor[1], s_7_38, c_8_39, c_7_7);
    divider_cell cell_8_39(s_8_39, c_8_39, divisor[0], dividend[23], c_7_7, c_7_7);
    assign div_result[23] = c_8_8;
    wire c_9_9, c_9_10, c_9_11, c_9_12, c_9_13, c_9_14, c_9_15, c_9_16, c_9_17, c_9_18, c_9_19, c_9_20, c_9_21, c_9_22, c_9_23, c_9_24, c_9_25, c_9_26, c_9_27, c_9_28, c_9_29, c_9_30, c_9_31, c_9_32, c_9_33, c_9_34, c_9_35, c_9_36, c_9_37, c_9_38, c_9_39, c_9_40;
    wire empty9, s_9_10, s_9_11, s_9_12, s_9_13, s_9_14, s_9_15, s_9_16, s_9_17, s_9_18, s_9_19, s_9_20, s_9_21, s_9_22, s_9_23, s_9_24, s_9_25, s_9_26, s_9_27, s_9_28, s_9_29, s_9_30, s_9_31, s_9_32, s_9_33, s_9_34, s_9_35, s_9_36, s_9_37, s_9_38, s_9_39, s_9_40;
    divider_cell cell_9_9(empty9, c_9_9, divisor[31], s_8_9, c_9_10, c_8_8);
    divider_cell cell_9_10(s_9_10, c_9_10, divisor[30], s_8_10, c_9_11, c_8_8);
    divider_cell cell_9_11(s_9_11, c_9_11, divisor[29], s_8_11, c_9_12, c_8_8);
    divider_cell cell_9_12(s_9_12, c_9_12, divisor[28], s_8_12, c_9_13, c_8_8);
    divider_cell cell_9_13(s_9_13, c_9_13, divisor[27], s_8_13, c_9_14, c_8_8);
    divider_cell cell_9_14(s_9_14, c_9_14, divisor[26], s_8_14, c_9_15, c_8_8);
    divider_cell cell_9_15(s_9_15, c_9_15, divisor[25], s_8_15, c_9_16, c_8_8);
    divider_cell cell_9_16(s_9_16, c_9_16, divisor[24], s_8_16, c_9_17, c_8_8);
    divider_cell cell_9_17(s_9_17, c_9_17, divisor[23], s_8_17, c_9_18, c_8_8);
    divider_cell cell_9_18(s_9_18, c_9_18, divisor[22], s_8_18, c_9_19, c_8_8);
    divider_cell cell_9_19(s_9_19, c_9_19, divisor[21], s_8_19, c_9_20, c_8_8);
    divider_cell cell_9_20(s_9_20, c_9_20, divisor[20], s_8_20, c_9_21, c_8_8);
    divider_cell cell_9_21(s_9_21, c_9_21, divisor[19], s_8_21, c_9_22, c_8_8);
    divider_cell cell_9_22(s_9_22, c_9_22, divisor[18], s_8_22, c_9_23, c_8_8);
    divider_cell cell_9_23(s_9_23, c_9_23, divisor[17], s_8_23, c_9_24, c_8_8);
    divider_cell cell_9_24(s_9_24, c_9_24, divisor[16], s_8_24, c_9_25, c_8_8);
    divider_cell cell_9_25(s_9_25, c_9_25, divisor[15], s_8_25, c_9_26, c_8_8);
    divider_cell cell_9_26(s_9_26, c_9_26, divisor[14], s_8_26, c_9_27, c_8_8);
    divider_cell cell_9_27(s_9_27, c_9_27, divisor[13], s_8_27, c_9_28, c_8_8);
    divider_cell cell_9_28(s_9_28, c_9_28, divisor[12], s_8_28, c_9_29, c_8_8);
    divider_cell cell_9_29(s_9_29, c_9_29, divisor[11], s_8_29, c_9_30, c_8_8);
    divider_cell cell_9_30(s_9_30, c_9_30, divisor[10], s_8_30, c_9_31, c_8_8);
    divider_cell cell_9_31(s_9_31, c_9_31, divisor[9], s_8_31, c_9_32, c_8_8);
    divider_cell cell_9_32(s_9_32, c_9_32, divisor[8], s_8_32, c_9_33, c_8_8);
    divider_cell cell_9_33(s_9_33, c_9_33, divisor[7], s_8_33, c_9_34, c_8_8);
    divider_cell cell_9_34(s_9_34, c_9_34, divisor[6], s_8_34, c_9_35, c_8_8);
    divider_cell cell_9_35(s_9_35, c_9_35, divisor[5], s_8_35, c_9_36, c_8_8);
    divider_cell cell_9_36(s_9_36, c_9_36, divisor[4], s_8_36, c_9_37, c_8_8);
    divider_cell cell_9_37(s_9_37, c_9_37, divisor[3], s_8_37, c_9_38, c_8_8);
    divider_cell cell_9_38(s_9_38, c_9_38, divisor[2], s_8_38, c_9_39, c_8_8);
    divider_cell cell_9_39(s_9_39, c_9_39, divisor[1], s_8_39, c_9_40, c_8_8);
    divider_cell cell_9_40(s_9_40, c_9_40, divisor[0], dividend[22], c_8_8, c_8_8);
    assign div_result[22] = c_9_9;
    wire c_10_10, c_10_11, c_10_12, c_10_13, c_10_14, c_10_15, c_10_16, c_10_17, c_10_18, c_10_19, c_10_20, c_10_21, c_10_22, c_10_23, c_10_24, c_10_25, c_10_26, c_10_27, c_10_28, c_10_29, c_10_30, c_10_31, c_10_32, c_10_33, c_10_34, c_10_35, c_10_36, c_10_37, c_10_38, c_10_39, c_10_40, c_10_41;
    wire empty10, s_10_11, s_10_12, s_10_13, s_10_14, s_10_15, s_10_16, s_10_17, s_10_18, s_10_19, s_10_20, s_10_21, s_10_22, s_10_23, s_10_24, s_10_25, s_10_26, s_10_27, s_10_28, s_10_29, s_10_30, s_10_31, s_10_32, s_10_33, s_10_34, s_10_35, s_10_36, s_10_37, s_10_38, s_10_39, s_10_40, s_10_41;
    divider_cell cell_10_10(empty10, c_10_10, divisor[31], s_9_10, c_10_11, c_9_9);
    divider_cell cell_10_11(s_10_11, c_10_11, divisor[30], s_9_11, c_10_12, c_9_9);
    divider_cell cell_10_12(s_10_12, c_10_12, divisor[29], s_9_12, c_10_13, c_9_9);
    divider_cell cell_10_13(s_10_13, c_10_13, divisor[28], s_9_13, c_10_14, c_9_9);
    divider_cell cell_10_14(s_10_14, c_10_14, divisor[27], s_9_14, c_10_15, c_9_9);
    divider_cell cell_10_15(s_10_15, c_10_15, divisor[26], s_9_15, c_10_16, c_9_9);
    divider_cell cell_10_16(s_10_16, c_10_16, divisor[25], s_9_16, c_10_17, c_9_9);
    divider_cell cell_10_17(s_10_17, c_10_17, divisor[24], s_9_17, c_10_18, c_9_9);
    divider_cell cell_10_18(s_10_18, c_10_18, divisor[23], s_9_18, c_10_19, c_9_9);
    divider_cell cell_10_19(s_10_19, c_10_19, divisor[22], s_9_19, c_10_20, c_9_9);
    divider_cell cell_10_20(s_10_20, c_10_20, divisor[21], s_9_20, c_10_21, c_9_9);
    divider_cell cell_10_21(s_10_21, c_10_21, divisor[20], s_9_21, c_10_22, c_9_9);
    divider_cell cell_10_22(s_10_22, c_10_22, divisor[19], s_9_22, c_10_23, c_9_9);
    divider_cell cell_10_23(s_10_23, c_10_23, divisor[18], s_9_23, c_10_24, c_9_9);
    divider_cell cell_10_24(s_10_24, c_10_24, divisor[17], s_9_24, c_10_25, c_9_9);
    divider_cell cell_10_25(s_10_25, c_10_25, divisor[16], s_9_25, c_10_26, c_9_9);
    divider_cell cell_10_26(s_10_26, c_10_26, divisor[15], s_9_26, c_10_27, c_9_9);
    divider_cell cell_10_27(s_10_27, c_10_27, divisor[14], s_9_27, c_10_28, c_9_9);
    divider_cell cell_10_28(s_10_28, c_10_28, divisor[13], s_9_28, c_10_29, c_9_9);
    divider_cell cell_10_29(s_10_29, c_10_29, divisor[12], s_9_29, c_10_30, c_9_9);
    divider_cell cell_10_30(s_10_30, c_10_30, divisor[11], s_9_30, c_10_31, c_9_9);
    divider_cell cell_10_31(s_10_31, c_10_31, divisor[10], s_9_31, c_10_32, c_9_9);
    divider_cell cell_10_32(s_10_32, c_10_32, divisor[9], s_9_32, c_10_33, c_9_9);
    divider_cell cell_10_33(s_10_33, c_10_33, divisor[8], s_9_33, c_10_34, c_9_9);
    divider_cell cell_10_34(s_10_34, c_10_34, divisor[7], s_9_34, c_10_35, c_9_9);
    divider_cell cell_10_35(s_10_35, c_10_35, divisor[6], s_9_35, c_10_36, c_9_9);
    divider_cell cell_10_36(s_10_36, c_10_36, divisor[5], s_9_36, c_10_37, c_9_9);
    divider_cell cell_10_37(s_10_37, c_10_37, divisor[4], s_9_37, c_10_38, c_9_9);
    divider_cell cell_10_38(s_10_38, c_10_38, divisor[3], s_9_38, c_10_39, c_9_9);
    divider_cell cell_10_39(s_10_39, c_10_39, divisor[2], s_9_39, c_10_40, c_9_9);
    divider_cell cell_10_40(s_10_40, c_10_40, divisor[1], s_9_40, c_10_41, c_9_9);
    divider_cell cell_10_41(s_10_41, c_10_41, divisor[0], dividend[21], c_9_9, c_9_9);
    assign div_result[21] = c_10_10;
    wire c_11_11, c_11_12, c_11_13, c_11_14, c_11_15, c_11_16, c_11_17, c_11_18, c_11_19, c_11_20, c_11_21, c_11_22, c_11_23, c_11_24, c_11_25, c_11_26, c_11_27, c_11_28, c_11_29, c_11_30, c_11_31, c_11_32, c_11_33, c_11_34, c_11_35, c_11_36, c_11_37, c_11_38, c_11_39, c_11_40, c_11_41, c_11_42;
    wire empty11, s_11_12, s_11_13, s_11_14, s_11_15, s_11_16, s_11_17, s_11_18, s_11_19, s_11_20, s_11_21, s_11_22, s_11_23, s_11_24, s_11_25, s_11_26, s_11_27, s_11_28, s_11_29, s_11_30, s_11_31, s_11_32, s_11_33, s_11_34, s_11_35, s_11_36, s_11_37, s_11_38, s_11_39, s_11_40, s_11_41, s_11_42;
    divider_cell cell_11_11(empty11, c_11_11, divisor[31], s_10_11, c_11_12, c_10_10);
    divider_cell cell_11_12(s_11_12, c_11_12, divisor[30], s_10_12, c_11_13, c_10_10);
    divider_cell cell_11_13(s_11_13, c_11_13, divisor[29], s_10_13, c_11_14, c_10_10);
    divider_cell cell_11_14(s_11_14, c_11_14, divisor[28], s_10_14, c_11_15, c_10_10);
    divider_cell cell_11_15(s_11_15, c_11_15, divisor[27], s_10_15, c_11_16, c_10_10);
    divider_cell cell_11_16(s_11_16, c_11_16, divisor[26], s_10_16, c_11_17, c_10_10);
    divider_cell cell_11_17(s_11_17, c_11_17, divisor[25], s_10_17, c_11_18, c_10_10);
    divider_cell cell_11_18(s_11_18, c_11_18, divisor[24], s_10_18, c_11_19, c_10_10);
    divider_cell cell_11_19(s_11_19, c_11_19, divisor[23], s_10_19, c_11_20, c_10_10);
    divider_cell cell_11_20(s_11_20, c_11_20, divisor[22], s_10_20, c_11_21, c_10_10);
    divider_cell cell_11_21(s_11_21, c_11_21, divisor[21], s_10_21, c_11_22, c_10_10);
    divider_cell cell_11_22(s_11_22, c_11_22, divisor[20], s_10_22, c_11_23, c_10_10);
    divider_cell cell_11_23(s_11_23, c_11_23, divisor[19], s_10_23, c_11_24, c_10_10);
    divider_cell cell_11_24(s_11_24, c_11_24, divisor[18], s_10_24, c_11_25, c_10_10);
    divider_cell cell_11_25(s_11_25, c_11_25, divisor[17], s_10_25, c_11_26, c_10_10);
    divider_cell cell_11_26(s_11_26, c_11_26, divisor[16], s_10_26, c_11_27, c_10_10);
    divider_cell cell_11_27(s_11_27, c_11_27, divisor[15], s_10_27, c_11_28, c_10_10);
    divider_cell cell_11_28(s_11_28, c_11_28, divisor[14], s_10_28, c_11_29, c_10_10);
    divider_cell cell_11_29(s_11_29, c_11_29, divisor[13], s_10_29, c_11_30, c_10_10);
    divider_cell cell_11_30(s_11_30, c_11_30, divisor[12], s_10_30, c_11_31, c_10_10);
    divider_cell cell_11_31(s_11_31, c_11_31, divisor[11], s_10_31, c_11_32, c_10_10);
    divider_cell cell_11_32(s_11_32, c_11_32, divisor[10], s_10_32, c_11_33, c_10_10);
    divider_cell cell_11_33(s_11_33, c_11_33, divisor[9], s_10_33, c_11_34, c_10_10);
    divider_cell cell_11_34(s_11_34, c_11_34, divisor[8], s_10_34, c_11_35, c_10_10);
    divider_cell cell_11_35(s_11_35, c_11_35, divisor[7], s_10_35, c_11_36, c_10_10);
    divider_cell cell_11_36(s_11_36, c_11_36, divisor[6], s_10_36, c_11_37, c_10_10);
    divider_cell cell_11_37(s_11_37, c_11_37, divisor[5], s_10_37, c_11_38, c_10_10);
    divider_cell cell_11_38(s_11_38, c_11_38, divisor[4], s_10_38, c_11_39, c_10_10);
    divider_cell cell_11_39(s_11_39, c_11_39, divisor[3], s_10_39, c_11_40, c_10_10);
    divider_cell cell_11_40(s_11_40, c_11_40, divisor[2], s_10_40, c_11_41, c_10_10);
    divider_cell cell_11_41(s_11_41, c_11_41, divisor[1], s_10_41, c_11_42, c_10_10);
    divider_cell cell_11_42(s_11_42, c_11_42, divisor[0], dividend[20], c_10_10, c_10_10);
    assign div_result[20] = c_11_11;
    wire c_12_12, c_12_13, c_12_14, c_12_15, c_12_16, c_12_17, c_12_18, c_12_19, c_12_20, c_12_21, c_12_22, c_12_23, c_12_24, c_12_25, c_12_26, c_12_27, c_12_28, c_12_29, c_12_30, c_12_31, c_12_32, c_12_33, c_12_34, c_12_35, c_12_36, c_12_37, c_12_38, c_12_39, c_12_40, c_12_41, c_12_42, c_12_43;
    wire empty12, s_12_13, s_12_14, s_12_15, s_12_16, s_12_17, s_12_18, s_12_19, s_12_20, s_12_21, s_12_22, s_12_23, s_12_24, s_12_25, s_12_26, s_12_27, s_12_28, s_12_29, s_12_30, s_12_31, s_12_32, s_12_33, s_12_34, s_12_35, s_12_36, s_12_37, s_12_38, s_12_39, s_12_40, s_12_41, s_12_42, s_12_43;
    divider_cell cell_12_12(empty12, c_12_12, divisor[31], s_11_12, c_12_13, c_11_11);
    divider_cell cell_12_13(s_12_13, c_12_13, divisor[30], s_11_13, c_12_14, c_11_11);
    divider_cell cell_12_14(s_12_14, c_12_14, divisor[29], s_11_14, c_12_15, c_11_11);
    divider_cell cell_12_15(s_12_15, c_12_15, divisor[28], s_11_15, c_12_16, c_11_11);
    divider_cell cell_12_16(s_12_16, c_12_16, divisor[27], s_11_16, c_12_17, c_11_11);
    divider_cell cell_12_17(s_12_17, c_12_17, divisor[26], s_11_17, c_12_18, c_11_11);
    divider_cell cell_12_18(s_12_18, c_12_18, divisor[25], s_11_18, c_12_19, c_11_11);
    divider_cell cell_12_19(s_12_19, c_12_19, divisor[24], s_11_19, c_12_20, c_11_11);
    divider_cell cell_12_20(s_12_20, c_12_20, divisor[23], s_11_20, c_12_21, c_11_11);
    divider_cell cell_12_21(s_12_21, c_12_21, divisor[22], s_11_21, c_12_22, c_11_11);
    divider_cell cell_12_22(s_12_22, c_12_22, divisor[21], s_11_22, c_12_23, c_11_11);
    divider_cell cell_12_23(s_12_23, c_12_23, divisor[20], s_11_23, c_12_24, c_11_11);
    divider_cell cell_12_24(s_12_24, c_12_24, divisor[19], s_11_24, c_12_25, c_11_11);
    divider_cell cell_12_25(s_12_25, c_12_25, divisor[18], s_11_25, c_12_26, c_11_11);
    divider_cell cell_12_26(s_12_26, c_12_26, divisor[17], s_11_26, c_12_27, c_11_11);
    divider_cell cell_12_27(s_12_27, c_12_27, divisor[16], s_11_27, c_12_28, c_11_11);
    divider_cell cell_12_28(s_12_28, c_12_28, divisor[15], s_11_28, c_12_29, c_11_11);
    divider_cell cell_12_29(s_12_29, c_12_29, divisor[14], s_11_29, c_12_30, c_11_11);
    divider_cell cell_12_30(s_12_30, c_12_30, divisor[13], s_11_30, c_12_31, c_11_11);
    divider_cell cell_12_31(s_12_31, c_12_31, divisor[12], s_11_31, c_12_32, c_11_11);
    divider_cell cell_12_32(s_12_32, c_12_32, divisor[11], s_11_32, c_12_33, c_11_11);
    divider_cell cell_12_33(s_12_33, c_12_33, divisor[10], s_11_33, c_12_34, c_11_11);
    divider_cell cell_12_34(s_12_34, c_12_34, divisor[9], s_11_34, c_12_35, c_11_11);
    divider_cell cell_12_35(s_12_35, c_12_35, divisor[8], s_11_35, c_12_36, c_11_11);
    divider_cell cell_12_36(s_12_36, c_12_36, divisor[7], s_11_36, c_12_37, c_11_11);
    divider_cell cell_12_37(s_12_37, c_12_37, divisor[6], s_11_37, c_12_38, c_11_11);
    divider_cell cell_12_38(s_12_38, c_12_38, divisor[5], s_11_38, c_12_39, c_11_11);
    divider_cell cell_12_39(s_12_39, c_12_39, divisor[4], s_11_39, c_12_40, c_11_11);
    divider_cell cell_12_40(s_12_40, c_12_40, divisor[3], s_11_40, c_12_41, c_11_11);
    divider_cell cell_12_41(s_12_41, c_12_41, divisor[2], s_11_41, c_12_42, c_11_11);
    divider_cell cell_12_42(s_12_42, c_12_42, divisor[1], s_11_42, c_12_43, c_11_11);
    divider_cell cell_12_43(s_12_43, c_12_43, divisor[0], dividend[19], c_11_11, c_11_11);
    assign div_result[19] = c_12_12;
    wire c_13_13, c_13_14, c_13_15, c_13_16, c_13_17, c_13_18, c_13_19, c_13_20, c_13_21, c_13_22, c_13_23, c_13_24, c_13_25, c_13_26, c_13_27, c_13_28, c_13_29, c_13_30, c_13_31, c_13_32, c_13_33, c_13_34, c_13_35, c_13_36, c_13_37, c_13_38, c_13_39, c_13_40, c_13_41, c_13_42, c_13_43, c_13_44;
    wire empty13, s_13_14, s_13_15, s_13_16, s_13_17, s_13_18, s_13_19, s_13_20, s_13_21, s_13_22, s_13_23, s_13_24, s_13_25, s_13_26, s_13_27, s_13_28, s_13_29, s_13_30, s_13_31, s_13_32, s_13_33, s_13_34, s_13_35, s_13_36, s_13_37, s_13_38, s_13_39, s_13_40, s_13_41, s_13_42, s_13_43, s_13_44;
    divider_cell cell_13_13(empty13, c_13_13, divisor[31], s_12_13, c_13_14, c_12_12);
    divider_cell cell_13_14(s_13_14, c_13_14, divisor[30], s_12_14, c_13_15, c_12_12);
    divider_cell cell_13_15(s_13_15, c_13_15, divisor[29], s_12_15, c_13_16, c_12_12);
    divider_cell cell_13_16(s_13_16, c_13_16, divisor[28], s_12_16, c_13_17, c_12_12);
    divider_cell cell_13_17(s_13_17, c_13_17, divisor[27], s_12_17, c_13_18, c_12_12);
    divider_cell cell_13_18(s_13_18, c_13_18, divisor[26], s_12_18, c_13_19, c_12_12);
    divider_cell cell_13_19(s_13_19, c_13_19, divisor[25], s_12_19, c_13_20, c_12_12);
    divider_cell cell_13_20(s_13_20, c_13_20, divisor[24], s_12_20, c_13_21, c_12_12);
    divider_cell cell_13_21(s_13_21, c_13_21, divisor[23], s_12_21, c_13_22, c_12_12);
    divider_cell cell_13_22(s_13_22, c_13_22, divisor[22], s_12_22, c_13_23, c_12_12);
    divider_cell cell_13_23(s_13_23, c_13_23, divisor[21], s_12_23, c_13_24, c_12_12);
    divider_cell cell_13_24(s_13_24, c_13_24, divisor[20], s_12_24, c_13_25, c_12_12);
    divider_cell cell_13_25(s_13_25, c_13_25, divisor[19], s_12_25, c_13_26, c_12_12);
    divider_cell cell_13_26(s_13_26, c_13_26, divisor[18], s_12_26, c_13_27, c_12_12);
    divider_cell cell_13_27(s_13_27, c_13_27, divisor[17], s_12_27, c_13_28, c_12_12);
    divider_cell cell_13_28(s_13_28, c_13_28, divisor[16], s_12_28, c_13_29, c_12_12);
    divider_cell cell_13_29(s_13_29, c_13_29, divisor[15], s_12_29, c_13_30, c_12_12);
    divider_cell cell_13_30(s_13_30, c_13_30, divisor[14], s_12_30, c_13_31, c_12_12);
    divider_cell cell_13_31(s_13_31, c_13_31, divisor[13], s_12_31, c_13_32, c_12_12);
    divider_cell cell_13_32(s_13_32, c_13_32, divisor[12], s_12_32, c_13_33, c_12_12);
    divider_cell cell_13_33(s_13_33, c_13_33, divisor[11], s_12_33, c_13_34, c_12_12);
    divider_cell cell_13_34(s_13_34, c_13_34, divisor[10], s_12_34, c_13_35, c_12_12);
    divider_cell cell_13_35(s_13_35, c_13_35, divisor[9], s_12_35, c_13_36, c_12_12);
    divider_cell cell_13_36(s_13_36, c_13_36, divisor[8], s_12_36, c_13_37, c_12_12);
    divider_cell cell_13_37(s_13_37, c_13_37, divisor[7], s_12_37, c_13_38, c_12_12);
    divider_cell cell_13_38(s_13_38, c_13_38, divisor[6], s_12_38, c_13_39, c_12_12);
    divider_cell cell_13_39(s_13_39, c_13_39, divisor[5], s_12_39, c_13_40, c_12_12);
    divider_cell cell_13_40(s_13_40, c_13_40, divisor[4], s_12_40, c_13_41, c_12_12);
    divider_cell cell_13_41(s_13_41, c_13_41, divisor[3], s_12_41, c_13_42, c_12_12);
    divider_cell cell_13_42(s_13_42, c_13_42, divisor[2], s_12_42, c_13_43, c_12_12);
    divider_cell cell_13_43(s_13_43, c_13_43, divisor[1], s_12_43, c_13_44, c_12_12);
    divider_cell cell_13_44(s_13_44, c_13_44, divisor[0], dividend[18], c_12_12, c_12_12);
    assign div_result[18] = c_13_13;
    wire c_14_14, c_14_15, c_14_16, c_14_17, c_14_18, c_14_19, c_14_20, c_14_21, c_14_22, c_14_23, c_14_24, c_14_25, c_14_26, c_14_27, c_14_28, c_14_29, c_14_30, c_14_31, c_14_32, c_14_33, c_14_34, c_14_35, c_14_36, c_14_37, c_14_38, c_14_39, c_14_40, c_14_41, c_14_42, c_14_43, c_14_44, c_14_45;
    wire empty14, s_14_15, s_14_16, s_14_17, s_14_18, s_14_19, s_14_20, s_14_21, s_14_22, s_14_23, s_14_24, s_14_25, s_14_26, s_14_27, s_14_28, s_14_29, s_14_30, s_14_31, s_14_32, s_14_33, s_14_34, s_14_35, s_14_36, s_14_37, s_14_38, s_14_39, s_14_40, s_14_41, s_14_42, s_14_43, s_14_44, s_14_45;
    divider_cell cell_14_14(empty14, c_14_14, divisor[31], s_13_14, c_14_15, c_13_13);
    divider_cell cell_14_15(s_14_15, c_14_15, divisor[30], s_13_15, c_14_16, c_13_13);
    divider_cell cell_14_16(s_14_16, c_14_16, divisor[29], s_13_16, c_14_17, c_13_13);
    divider_cell cell_14_17(s_14_17, c_14_17, divisor[28], s_13_17, c_14_18, c_13_13);
    divider_cell cell_14_18(s_14_18, c_14_18, divisor[27], s_13_18, c_14_19, c_13_13);
    divider_cell cell_14_19(s_14_19, c_14_19, divisor[26], s_13_19, c_14_20, c_13_13);
    divider_cell cell_14_20(s_14_20, c_14_20, divisor[25], s_13_20, c_14_21, c_13_13);
    divider_cell cell_14_21(s_14_21, c_14_21, divisor[24], s_13_21, c_14_22, c_13_13);
    divider_cell cell_14_22(s_14_22, c_14_22, divisor[23], s_13_22, c_14_23, c_13_13);
    divider_cell cell_14_23(s_14_23, c_14_23, divisor[22], s_13_23, c_14_24, c_13_13);
    divider_cell cell_14_24(s_14_24, c_14_24, divisor[21], s_13_24, c_14_25, c_13_13);
    divider_cell cell_14_25(s_14_25, c_14_25, divisor[20], s_13_25, c_14_26, c_13_13);
    divider_cell cell_14_26(s_14_26, c_14_26, divisor[19], s_13_26, c_14_27, c_13_13);
    divider_cell cell_14_27(s_14_27, c_14_27, divisor[18], s_13_27, c_14_28, c_13_13);
    divider_cell cell_14_28(s_14_28, c_14_28, divisor[17], s_13_28, c_14_29, c_13_13);
    divider_cell cell_14_29(s_14_29, c_14_29, divisor[16], s_13_29, c_14_30, c_13_13);
    divider_cell cell_14_30(s_14_30, c_14_30, divisor[15], s_13_30, c_14_31, c_13_13);
    divider_cell cell_14_31(s_14_31, c_14_31, divisor[14], s_13_31, c_14_32, c_13_13);
    divider_cell cell_14_32(s_14_32, c_14_32, divisor[13], s_13_32, c_14_33, c_13_13);
    divider_cell cell_14_33(s_14_33, c_14_33, divisor[12], s_13_33, c_14_34, c_13_13);
    divider_cell cell_14_34(s_14_34, c_14_34, divisor[11], s_13_34, c_14_35, c_13_13);
    divider_cell cell_14_35(s_14_35, c_14_35, divisor[10], s_13_35, c_14_36, c_13_13);
    divider_cell cell_14_36(s_14_36, c_14_36, divisor[9], s_13_36, c_14_37, c_13_13);
    divider_cell cell_14_37(s_14_37, c_14_37, divisor[8], s_13_37, c_14_38, c_13_13);
    divider_cell cell_14_38(s_14_38, c_14_38, divisor[7], s_13_38, c_14_39, c_13_13);
    divider_cell cell_14_39(s_14_39, c_14_39, divisor[6], s_13_39, c_14_40, c_13_13);
    divider_cell cell_14_40(s_14_40, c_14_40, divisor[5], s_13_40, c_14_41, c_13_13);
    divider_cell cell_14_41(s_14_41, c_14_41, divisor[4], s_13_41, c_14_42, c_13_13);
    divider_cell cell_14_42(s_14_42, c_14_42, divisor[3], s_13_42, c_14_43, c_13_13);
    divider_cell cell_14_43(s_14_43, c_14_43, divisor[2], s_13_43, c_14_44, c_13_13);
    divider_cell cell_14_44(s_14_44, c_14_44, divisor[1], s_13_44, c_14_45, c_13_13);
    divider_cell cell_14_45(s_14_45, c_14_45, divisor[0], dividend[17], c_13_13, c_13_13);
    assign div_result[17] = c_14_14;
    wire c_15_15, c_15_16, c_15_17, c_15_18, c_15_19, c_15_20, c_15_21, c_15_22, c_15_23, c_15_24, c_15_25, c_15_26, c_15_27, c_15_28, c_15_29, c_15_30, c_15_31, c_15_32, c_15_33, c_15_34, c_15_35, c_15_36, c_15_37, c_15_38, c_15_39, c_15_40, c_15_41, c_15_42, c_15_43, c_15_44, c_15_45, c_15_46;
    wire empty15, s_15_16, s_15_17, s_15_18, s_15_19, s_15_20, s_15_21, s_15_22, s_15_23, s_15_24, s_15_25, s_15_26, s_15_27, s_15_28, s_15_29, s_15_30, s_15_31, s_15_32, s_15_33, s_15_34, s_15_35, s_15_36, s_15_37, s_15_38, s_15_39, s_15_40, s_15_41, s_15_42, s_15_43, s_15_44, s_15_45, s_15_46;
    divider_cell cell_15_15(empty15, c_15_15, divisor[31], s_14_15, c_15_16, c_14_14);
    divider_cell cell_15_16(s_15_16, c_15_16, divisor[30], s_14_16, c_15_17, c_14_14);
    divider_cell cell_15_17(s_15_17, c_15_17, divisor[29], s_14_17, c_15_18, c_14_14);
    divider_cell cell_15_18(s_15_18, c_15_18, divisor[28], s_14_18, c_15_19, c_14_14);
    divider_cell cell_15_19(s_15_19, c_15_19, divisor[27], s_14_19, c_15_20, c_14_14);
    divider_cell cell_15_20(s_15_20, c_15_20, divisor[26], s_14_20, c_15_21, c_14_14);
    divider_cell cell_15_21(s_15_21, c_15_21, divisor[25], s_14_21, c_15_22, c_14_14);
    divider_cell cell_15_22(s_15_22, c_15_22, divisor[24], s_14_22, c_15_23, c_14_14);
    divider_cell cell_15_23(s_15_23, c_15_23, divisor[23], s_14_23, c_15_24, c_14_14);
    divider_cell cell_15_24(s_15_24, c_15_24, divisor[22], s_14_24, c_15_25, c_14_14);
    divider_cell cell_15_25(s_15_25, c_15_25, divisor[21], s_14_25, c_15_26, c_14_14);
    divider_cell cell_15_26(s_15_26, c_15_26, divisor[20], s_14_26, c_15_27, c_14_14);
    divider_cell cell_15_27(s_15_27, c_15_27, divisor[19], s_14_27, c_15_28, c_14_14);
    divider_cell cell_15_28(s_15_28, c_15_28, divisor[18], s_14_28, c_15_29, c_14_14);
    divider_cell cell_15_29(s_15_29, c_15_29, divisor[17], s_14_29, c_15_30, c_14_14);
    divider_cell cell_15_30(s_15_30, c_15_30, divisor[16], s_14_30, c_15_31, c_14_14);
    divider_cell cell_15_31(s_15_31, c_15_31, divisor[15], s_14_31, c_15_32, c_14_14);
    divider_cell cell_15_32(s_15_32, c_15_32, divisor[14], s_14_32, c_15_33, c_14_14);
    divider_cell cell_15_33(s_15_33, c_15_33, divisor[13], s_14_33, c_15_34, c_14_14);
    divider_cell cell_15_34(s_15_34, c_15_34, divisor[12], s_14_34, c_15_35, c_14_14);
    divider_cell cell_15_35(s_15_35, c_15_35, divisor[11], s_14_35, c_15_36, c_14_14);
    divider_cell cell_15_36(s_15_36, c_15_36, divisor[10], s_14_36, c_15_37, c_14_14);
    divider_cell cell_15_37(s_15_37, c_15_37, divisor[9], s_14_37, c_15_38, c_14_14);
    divider_cell cell_15_38(s_15_38, c_15_38, divisor[8], s_14_38, c_15_39, c_14_14);
    divider_cell cell_15_39(s_15_39, c_15_39, divisor[7], s_14_39, c_15_40, c_14_14);
    divider_cell cell_15_40(s_15_40, c_15_40, divisor[6], s_14_40, c_15_41, c_14_14);
    divider_cell cell_15_41(s_15_41, c_15_41, divisor[5], s_14_41, c_15_42, c_14_14);
    divider_cell cell_15_42(s_15_42, c_15_42, divisor[4], s_14_42, c_15_43, c_14_14);
    divider_cell cell_15_43(s_15_43, c_15_43, divisor[3], s_14_43, c_15_44, c_14_14);
    divider_cell cell_15_44(s_15_44, c_15_44, divisor[2], s_14_44, c_15_45, c_14_14);
    divider_cell cell_15_45(s_15_45, c_15_45, divisor[1], s_14_45, c_15_46, c_14_14);
    divider_cell cell_15_46(s_15_46, c_15_46, divisor[0], dividend[16], c_14_14, c_14_14);
    assign div_result[16] = c_15_15;
    wire c_16_16, c_16_17, c_16_18, c_16_19, c_16_20, c_16_21, c_16_22, c_16_23, c_16_24, c_16_25, c_16_26, c_16_27, c_16_28, c_16_29, c_16_30, c_16_31, c_16_32, c_16_33, c_16_34, c_16_35, c_16_36, c_16_37, c_16_38, c_16_39, c_16_40, c_16_41, c_16_42, c_16_43, c_16_44, c_16_45, c_16_46, c_16_47;
    wire empty16, s_16_17, s_16_18, s_16_19, s_16_20, s_16_21, s_16_22, s_16_23, s_16_24, s_16_25, s_16_26, s_16_27, s_16_28, s_16_29, s_16_30, s_16_31, s_16_32, s_16_33, s_16_34, s_16_35, s_16_36, s_16_37, s_16_38, s_16_39, s_16_40, s_16_41, s_16_42, s_16_43, s_16_44, s_16_45, s_16_46, s_16_47;
    divider_cell cell_16_16(empty16, c_16_16, divisor[31], s_15_16, c_16_17, c_15_15);
    divider_cell cell_16_17(s_16_17, c_16_17, divisor[30], s_15_17, c_16_18, c_15_15);
    divider_cell cell_16_18(s_16_18, c_16_18, divisor[29], s_15_18, c_16_19, c_15_15);
    divider_cell cell_16_19(s_16_19, c_16_19, divisor[28], s_15_19, c_16_20, c_15_15);
    divider_cell cell_16_20(s_16_20, c_16_20, divisor[27], s_15_20, c_16_21, c_15_15);
    divider_cell cell_16_21(s_16_21, c_16_21, divisor[26], s_15_21, c_16_22, c_15_15);
    divider_cell cell_16_22(s_16_22, c_16_22, divisor[25], s_15_22, c_16_23, c_15_15);
    divider_cell cell_16_23(s_16_23, c_16_23, divisor[24], s_15_23, c_16_24, c_15_15);
    divider_cell cell_16_24(s_16_24, c_16_24, divisor[23], s_15_24, c_16_25, c_15_15);
    divider_cell cell_16_25(s_16_25, c_16_25, divisor[22], s_15_25, c_16_26, c_15_15);
    divider_cell cell_16_26(s_16_26, c_16_26, divisor[21], s_15_26, c_16_27, c_15_15);
    divider_cell cell_16_27(s_16_27, c_16_27, divisor[20], s_15_27, c_16_28, c_15_15);
    divider_cell cell_16_28(s_16_28, c_16_28, divisor[19], s_15_28, c_16_29, c_15_15);
    divider_cell cell_16_29(s_16_29, c_16_29, divisor[18], s_15_29, c_16_30, c_15_15);
    divider_cell cell_16_30(s_16_30, c_16_30, divisor[17], s_15_30, c_16_31, c_15_15);
    divider_cell cell_16_31(s_16_31, c_16_31, divisor[16], s_15_31, c_16_32, c_15_15);
    divider_cell cell_16_32(s_16_32, c_16_32, divisor[15], s_15_32, c_16_33, c_15_15);
    divider_cell cell_16_33(s_16_33, c_16_33, divisor[14], s_15_33, c_16_34, c_15_15);
    divider_cell cell_16_34(s_16_34, c_16_34, divisor[13], s_15_34, c_16_35, c_15_15);
    divider_cell cell_16_35(s_16_35, c_16_35, divisor[12], s_15_35, c_16_36, c_15_15);
    divider_cell cell_16_36(s_16_36, c_16_36, divisor[11], s_15_36, c_16_37, c_15_15);
    divider_cell cell_16_37(s_16_37, c_16_37, divisor[10], s_15_37, c_16_38, c_15_15);
    divider_cell cell_16_38(s_16_38, c_16_38, divisor[9], s_15_38, c_16_39, c_15_15);
    divider_cell cell_16_39(s_16_39, c_16_39, divisor[8], s_15_39, c_16_40, c_15_15);
    divider_cell cell_16_40(s_16_40, c_16_40, divisor[7], s_15_40, c_16_41, c_15_15);
    divider_cell cell_16_41(s_16_41, c_16_41, divisor[6], s_15_41, c_16_42, c_15_15);
    divider_cell cell_16_42(s_16_42, c_16_42, divisor[5], s_15_42, c_16_43, c_15_15);
    divider_cell cell_16_43(s_16_43, c_16_43, divisor[4], s_15_43, c_16_44, c_15_15);
    divider_cell cell_16_44(s_16_44, c_16_44, divisor[3], s_15_44, c_16_45, c_15_15);
    divider_cell cell_16_45(s_16_45, c_16_45, divisor[2], s_15_45, c_16_46, c_15_15);
    divider_cell cell_16_46(s_16_46, c_16_46, divisor[1], s_15_46, c_16_47, c_15_15);
    divider_cell cell_16_47(s_16_47, c_16_47, divisor[0], dividend[15], c_15_15, c_15_15);
    assign div_result[15] = c_16_16;
    wire c_17_17, c_17_18, c_17_19, c_17_20, c_17_21, c_17_22, c_17_23, c_17_24, c_17_25, c_17_26, c_17_27, c_17_28, c_17_29, c_17_30, c_17_31, c_17_32, c_17_33, c_17_34, c_17_35, c_17_36, c_17_37, c_17_38, c_17_39, c_17_40, c_17_41, c_17_42, c_17_43, c_17_44, c_17_45, c_17_46, c_17_47, c_17_48;
    wire empty17, s_17_18, s_17_19, s_17_20, s_17_21, s_17_22, s_17_23, s_17_24, s_17_25, s_17_26, s_17_27, s_17_28, s_17_29, s_17_30, s_17_31, s_17_32, s_17_33, s_17_34, s_17_35, s_17_36, s_17_37, s_17_38, s_17_39, s_17_40, s_17_41, s_17_42, s_17_43, s_17_44, s_17_45, s_17_46, s_17_47, s_17_48;
    divider_cell cell_17_17(empty17, c_17_17, divisor[31], s_16_17, c_17_18, c_16_16);
    divider_cell cell_17_18(s_17_18, c_17_18, divisor[30], s_16_18, c_17_19, c_16_16);
    divider_cell cell_17_19(s_17_19, c_17_19, divisor[29], s_16_19, c_17_20, c_16_16);
    divider_cell cell_17_20(s_17_20, c_17_20, divisor[28], s_16_20, c_17_21, c_16_16);
    divider_cell cell_17_21(s_17_21, c_17_21, divisor[27], s_16_21, c_17_22, c_16_16);
    divider_cell cell_17_22(s_17_22, c_17_22, divisor[26], s_16_22, c_17_23, c_16_16);
    divider_cell cell_17_23(s_17_23, c_17_23, divisor[25], s_16_23, c_17_24, c_16_16);
    divider_cell cell_17_24(s_17_24, c_17_24, divisor[24], s_16_24, c_17_25, c_16_16);
    divider_cell cell_17_25(s_17_25, c_17_25, divisor[23], s_16_25, c_17_26, c_16_16);
    divider_cell cell_17_26(s_17_26, c_17_26, divisor[22], s_16_26, c_17_27, c_16_16);
    divider_cell cell_17_27(s_17_27, c_17_27, divisor[21], s_16_27, c_17_28, c_16_16);
    divider_cell cell_17_28(s_17_28, c_17_28, divisor[20], s_16_28, c_17_29, c_16_16);
    divider_cell cell_17_29(s_17_29, c_17_29, divisor[19], s_16_29, c_17_30, c_16_16);
    divider_cell cell_17_30(s_17_30, c_17_30, divisor[18], s_16_30, c_17_31, c_16_16);
    divider_cell cell_17_31(s_17_31, c_17_31, divisor[17], s_16_31, c_17_32, c_16_16);
    divider_cell cell_17_32(s_17_32, c_17_32, divisor[16], s_16_32, c_17_33, c_16_16);
    divider_cell cell_17_33(s_17_33, c_17_33, divisor[15], s_16_33, c_17_34, c_16_16);
    divider_cell cell_17_34(s_17_34, c_17_34, divisor[14], s_16_34, c_17_35, c_16_16);
    divider_cell cell_17_35(s_17_35, c_17_35, divisor[13], s_16_35, c_17_36, c_16_16);
    divider_cell cell_17_36(s_17_36, c_17_36, divisor[12], s_16_36, c_17_37, c_16_16);
    divider_cell cell_17_37(s_17_37, c_17_37, divisor[11], s_16_37, c_17_38, c_16_16);
    divider_cell cell_17_38(s_17_38, c_17_38, divisor[10], s_16_38, c_17_39, c_16_16);
    divider_cell cell_17_39(s_17_39, c_17_39, divisor[9], s_16_39, c_17_40, c_16_16);
    divider_cell cell_17_40(s_17_40, c_17_40, divisor[8], s_16_40, c_17_41, c_16_16);
    divider_cell cell_17_41(s_17_41, c_17_41, divisor[7], s_16_41, c_17_42, c_16_16);
    divider_cell cell_17_42(s_17_42, c_17_42, divisor[6], s_16_42, c_17_43, c_16_16);
    divider_cell cell_17_43(s_17_43, c_17_43, divisor[5], s_16_43, c_17_44, c_16_16);
    divider_cell cell_17_44(s_17_44, c_17_44, divisor[4], s_16_44, c_17_45, c_16_16);
    divider_cell cell_17_45(s_17_45, c_17_45, divisor[3], s_16_45, c_17_46, c_16_16);
    divider_cell cell_17_46(s_17_46, c_17_46, divisor[2], s_16_46, c_17_47, c_16_16);
    divider_cell cell_17_47(s_17_47, c_17_47, divisor[1], s_16_47, c_17_48, c_16_16);
    divider_cell cell_17_48(s_17_48, c_17_48, divisor[0], dividend[14], c_16_16, c_16_16);
    assign div_result[14] = c_17_17;
    wire c_18_18, c_18_19, c_18_20, c_18_21, c_18_22, c_18_23, c_18_24, c_18_25, c_18_26, c_18_27, c_18_28, c_18_29, c_18_30, c_18_31, c_18_32, c_18_33, c_18_34, c_18_35, c_18_36, c_18_37, c_18_38, c_18_39, c_18_40, c_18_41, c_18_42, c_18_43, c_18_44, c_18_45, c_18_46, c_18_47, c_18_48, c_18_49;
    wire empty18, s_18_19, s_18_20, s_18_21, s_18_22, s_18_23, s_18_24, s_18_25, s_18_26, s_18_27, s_18_28, s_18_29, s_18_30, s_18_31, s_18_32, s_18_33, s_18_34, s_18_35, s_18_36, s_18_37, s_18_38, s_18_39, s_18_40, s_18_41, s_18_42, s_18_43, s_18_44, s_18_45, s_18_46, s_18_47, s_18_48, s_18_49;
    divider_cell cell_18_18(empty18, c_18_18, divisor[31], s_17_18, c_18_19, c_17_17);
    divider_cell cell_18_19(s_18_19, c_18_19, divisor[30], s_17_19, c_18_20, c_17_17);
    divider_cell cell_18_20(s_18_20, c_18_20, divisor[29], s_17_20, c_18_21, c_17_17);
    divider_cell cell_18_21(s_18_21, c_18_21, divisor[28], s_17_21, c_18_22, c_17_17);
    divider_cell cell_18_22(s_18_22, c_18_22, divisor[27], s_17_22, c_18_23, c_17_17);
    divider_cell cell_18_23(s_18_23, c_18_23, divisor[26], s_17_23, c_18_24, c_17_17);
    divider_cell cell_18_24(s_18_24, c_18_24, divisor[25], s_17_24, c_18_25, c_17_17);
    divider_cell cell_18_25(s_18_25, c_18_25, divisor[24], s_17_25, c_18_26, c_17_17);
    divider_cell cell_18_26(s_18_26, c_18_26, divisor[23], s_17_26, c_18_27, c_17_17);
    divider_cell cell_18_27(s_18_27, c_18_27, divisor[22], s_17_27, c_18_28, c_17_17);
    divider_cell cell_18_28(s_18_28, c_18_28, divisor[21], s_17_28, c_18_29, c_17_17);
    divider_cell cell_18_29(s_18_29, c_18_29, divisor[20], s_17_29, c_18_30, c_17_17);
    divider_cell cell_18_30(s_18_30, c_18_30, divisor[19], s_17_30, c_18_31, c_17_17);
    divider_cell cell_18_31(s_18_31, c_18_31, divisor[18], s_17_31, c_18_32, c_17_17);
    divider_cell cell_18_32(s_18_32, c_18_32, divisor[17], s_17_32, c_18_33, c_17_17);
    divider_cell cell_18_33(s_18_33, c_18_33, divisor[16], s_17_33, c_18_34, c_17_17);
    divider_cell cell_18_34(s_18_34, c_18_34, divisor[15], s_17_34, c_18_35, c_17_17);
    divider_cell cell_18_35(s_18_35, c_18_35, divisor[14], s_17_35, c_18_36, c_17_17);
    divider_cell cell_18_36(s_18_36, c_18_36, divisor[13], s_17_36, c_18_37, c_17_17);
    divider_cell cell_18_37(s_18_37, c_18_37, divisor[12], s_17_37, c_18_38, c_17_17);
    divider_cell cell_18_38(s_18_38, c_18_38, divisor[11], s_17_38, c_18_39, c_17_17);
    divider_cell cell_18_39(s_18_39, c_18_39, divisor[10], s_17_39, c_18_40, c_17_17);
    divider_cell cell_18_40(s_18_40, c_18_40, divisor[9], s_17_40, c_18_41, c_17_17);
    divider_cell cell_18_41(s_18_41, c_18_41, divisor[8], s_17_41, c_18_42, c_17_17);
    divider_cell cell_18_42(s_18_42, c_18_42, divisor[7], s_17_42, c_18_43, c_17_17);
    divider_cell cell_18_43(s_18_43, c_18_43, divisor[6], s_17_43, c_18_44, c_17_17);
    divider_cell cell_18_44(s_18_44, c_18_44, divisor[5], s_17_44, c_18_45, c_17_17);
    divider_cell cell_18_45(s_18_45, c_18_45, divisor[4], s_17_45, c_18_46, c_17_17);
    divider_cell cell_18_46(s_18_46, c_18_46, divisor[3], s_17_46, c_18_47, c_17_17);
    divider_cell cell_18_47(s_18_47, c_18_47, divisor[2], s_17_47, c_18_48, c_17_17);
    divider_cell cell_18_48(s_18_48, c_18_48, divisor[1], s_17_48, c_18_49, c_17_17);
    divider_cell cell_18_49(s_18_49, c_18_49, divisor[0], dividend[13], c_17_17, c_17_17);
    assign div_result[13] = c_18_18;
    wire c_19_19, c_19_20, c_19_21, c_19_22, c_19_23, c_19_24, c_19_25, c_19_26, c_19_27, c_19_28, c_19_29, c_19_30, c_19_31, c_19_32, c_19_33, c_19_34, c_19_35, c_19_36, c_19_37, c_19_38, c_19_39, c_19_40, c_19_41, c_19_42, c_19_43, c_19_44, c_19_45, c_19_46, c_19_47, c_19_48, c_19_49, c_19_50;
    wire empty19, s_19_20, s_19_21, s_19_22, s_19_23, s_19_24, s_19_25, s_19_26, s_19_27, s_19_28, s_19_29, s_19_30, s_19_31, s_19_32, s_19_33, s_19_34, s_19_35, s_19_36, s_19_37, s_19_38, s_19_39, s_19_40, s_19_41, s_19_42, s_19_43, s_19_44, s_19_45, s_19_46, s_19_47, s_19_48, s_19_49, s_19_50;
    divider_cell cell_19_19(empty19, c_19_19, divisor[31], s_18_19, c_19_20, c_18_18);
    divider_cell cell_19_20(s_19_20, c_19_20, divisor[30], s_18_20, c_19_21, c_18_18);
    divider_cell cell_19_21(s_19_21, c_19_21, divisor[29], s_18_21, c_19_22, c_18_18);
    divider_cell cell_19_22(s_19_22, c_19_22, divisor[28], s_18_22, c_19_23, c_18_18);
    divider_cell cell_19_23(s_19_23, c_19_23, divisor[27], s_18_23, c_19_24, c_18_18);
    divider_cell cell_19_24(s_19_24, c_19_24, divisor[26], s_18_24, c_19_25, c_18_18);
    divider_cell cell_19_25(s_19_25, c_19_25, divisor[25], s_18_25, c_19_26, c_18_18);
    divider_cell cell_19_26(s_19_26, c_19_26, divisor[24], s_18_26, c_19_27, c_18_18);
    divider_cell cell_19_27(s_19_27, c_19_27, divisor[23], s_18_27, c_19_28, c_18_18);
    divider_cell cell_19_28(s_19_28, c_19_28, divisor[22], s_18_28, c_19_29, c_18_18);
    divider_cell cell_19_29(s_19_29, c_19_29, divisor[21], s_18_29, c_19_30, c_18_18);
    divider_cell cell_19_30(s_19_30, c_19_30, divisor[20], s_18_30, c_19_31, c_18_18);
    divider_cell cell_19_31(s_19_31, c_19_31, divisor[19], s_18_31, c_19_32, c_18_18);
    divider_cell cell_19_32(s_19_32, c_19_32, divisor[18], s_18_32, c_19_33, c_18_18);
    divider_cell cell_19_33(s_19_33, c_19_33, divisor[17], s_18_33, c_19_34, c_18_18);
    divider_cell cell_19_34(s_19_34, c_19_34, divisor[16], s_18_34, c_19_35, c_18_18);
    divider_cell cell_19_35(s_19_35, c_19_35, divisor[15], s_18_35, c_19_36, c_18_18);
    divider_cell cell_19_36(s_19_36, c_19_36, divisor[14], s_18_36, c_19_37, c_18_18);
    divider_cell cell_19_37(s_19_37, c_19_37, divisor[13], s_18_37, c_19_38, c_18_18);
    divider_cell cell_19_38(s_19_38, c_19_38, divisor[12], s_18_38, c_19_39, c_18_18);
    divider_cell cell_19_39(s_19_39, c_19_39, divisor[11], s_18_39, c_19_40, c_18_18);
    divider_cell cell_19_40(s_19_40, c_19_40, divisor[10], s_18_40, c_19_41, c_18_18);
    divider_cell cell_19_41(s_19_41, c_19_41, divisor[9], s_18_41, c_19_42, c_18_18);
    divider_cell cell_19_42(s_19_42, c_19_42, divisor[8], s_18_42, c_19_43, c_18_18);
    divider_cell cell_19_43(s_19_43, c_19_43, divisor[7], s_18_43, c_19_44, c_18_18);
    divider_cell cell_19_44(s_19_44, c_19_44, divisor[6], s_18_44, c_19_45, c_18_18);
    divider_cell cell_19_45(s_19_45, c_19_45, divisor[5], s_18_45, c_19_46, c_18_18);
    divider_cell cell_19_46(s_19_46, c_19_46, divisor[4], s_18_46, c_19_47, c_18_18);
    divider_cell cell_19_47(s_19_47, c_19_47, divisor[3], s_18_47, c_19_48, c_18_18);
    divider_cell cell_19_48(s_19_48, c_19_48, divisor[2], s_18_48, c_19_49, c_18_18);
    divider_cell cell_19_49(s_19_49, c_19_49, divisor[1], s_18_49, c_19_50, c_18_18);
    divider_cell cell_19_50(s_19_50, c_19_50, divisor[0], dividend[12], c_18_18, c_18_18);
    assign div_result[12] = c_19_19;
    wire c_20_20, c_20_21, c_20_22, c_20_23, c_20_24, c_20_25, c_20_26, c_20_27, c_20_28, c_20_29, c_20_30, c_20_31, c_20_32, c_20_33, c_20_34, c_20_35, c_20_36, c_20_37, c_20_38, c_20_39, c_20_40, c_20_41, c_20_42, c_20_43, c_20_44, c_20_45, c_20_46, c_20_47, c_20_48, c_20_49, c_20_50, c_20_51;
    wire empty20, s_20_21, s_20_22, s_20_23, s_20_24, s_20_25, s_20_26, s_20_27, s_20_28, s_20_29, s_20_30, s_20_31, s_20_32, s_20_33, s_20_34, s_20_35, s_20_36, s_20_37, s_20_38, s_20_39, s_20_40, s_20_41, s_20_42, s_20_43, s_20_44, s_20_45, s_20_46, s_20_47, s_20_48, s_20_49, s_20_50, s_20_51;
    divider_cell cell_20_20(empty20, c_20_20, divisor[31], s_19_20, c_20_21, c_19_19);
    divider_cell cell_20_21(s_20_21, c_20_21, divisor[30], s_19_21, c_20_22, c_19_19);
    divider_cell cell_20_22(s_20_22, c_20_22, divisor[29], s_19_22, c_20_23, c_19_19);
    divider_cell cell_20_23(s_20_23, c_20_23, divisor[28], s_19_23, c_20_24, c_19_19);
    divider_cell cell_20_24(s_20_24, c_20_24, divisor[27], s_19_24, c_20_25, c_19_19);
    divider_cell cell_20_25(s_20_25, c_20_25, divisor[26], s_19_25, c_20_26, c_19_19);
    divider_cell cell_20_26(s_20_26, c_20_26, divisor[25], s_19_26, c_20_27, c_19_19);
    divider_cell cell_20_27(s_20_27, c_20_27, divisor[24], s_19_27, c_20_28, c_19_19);
    divider_cell cell_20_28(s_20_28, c_20_28, divisor[23], s_19_28, c_20_29, c_19_19);
    divider_cell cell_20_29(s_20_29, c_20_29, divisor[22], s_19_29, c_20_30, c_19_19);
    divider_cell cell_20_30(s_20_30, c_20_30, divisor[21], s_19_30, c_20_31, c_19_19);
    divider_cell cell_20_31(s_20_31, c_20_31, divisor[20], s_19_31, c_20_32, c_19_19);
    divider_cell cell_20_32(s_20_32, c_20_32, divisor[19], s_19_32, c_20_33, c_19_19);
    divider_cell cell_20_33(s_20_33, c_20_33, divisor[18], s_19_33, c_20_34, c_19_19);
    divider_cell cell_20_34(s_20_34, c_20_34, divisor[17], s_19_34, c_20_35, c_19_19);
    divider_cell cell_20_35(s_20_35, c_20_35, divisor[16], s_19_35, c_20_36, c_19_19);
    divider_cell cell_20_36(s_20_36, c_20_36, divisor[15], s_19_36, c_20_37, c_19_19);
    divider_cell cell_20_37(s_20_37, c_20_37, divisor[14], s_19_37, c_20_38, c_19_19);
    divider_cell cell_20_38(s_20_38, c_20_38, divisor[13], s_19_38, c_20_39, c_19_19);
    divider_cell cell_20_39(s_20_39, c_20_39, divisor[12], s_19_39, c_20_40, c_19_19);
    divider_cell cell_20_40(s_20_40, c_20_40, divisor[11], s_19_40, c_20_41, c_19_19);
    divider_cell cell_20_41(s_20_41, c_20_41, divisor[10], s_19_41, c_20_42, c_19_19);
    divider_cell cell_20_42(s_20_42, c_20_42, divisor[9], s_19_42, c_20_43, c_19_19);
    divider_cell cell_20_43(s_20_43, c_20_43, divisor[8], s_19_43, c_20_44, c_19_19);
    divider_cell cell_20_44(s_20_44, c_20_44, divisor[7], s_19_44, c_20_45, c_19_19);
    divider_cell cell_20_45(s_20_45, c_20_45, divisor[6], s_19_45, c_20_46, c_19_19);
    divider_cell cell_20_46(s_20_46, c_20_46, divisor[5], s_19_46, c_20_47, c_19_19);
    divider_cell cell_20_47(s_20_47, c_20_47, divisor[4], s_19_47, c_20_48, c_19_19);
    divider_cell cell_20_48(s_20_48, c_20_48, divisor[3], s_19_48, c_20_49, c_19_19);
    divider_cell cell_20_49(s_20_49, c_20_49, divisor[2], s_19_49, c_20_50, c_19_19);
    divider_cell cell_20_50(s_20_50, c_20_50, divisor[1], s_19_50, c_20_51, c_19_19);
    divider_cell cell_20_51(s_20_51, c_20_51, divisor[0], dividend[11], c_19_19, c_19_19);
    assign div_result[11] = c_20_20;
    wire c_21_21, c_21_22, c_21_23, c_21_24, c_21_25, c_21_26, c_21_27, c_21_28, c_21_29, c_21_30, c_21_31, c_21_32, c_21_33, c_21_34, c_21_35, c_21_36, c_21_37, c_21_38, c_21_39, c_21_40, c_21_41, c_21_42, c_21_43, c_21_44, c_21_45, c_21_46, c_21_47, c_21_48, c_21_49, c_21_50, c_21_51, c_21_52;
    wire empty21, s_21_22, s_21_23, s_21_24, s_21_25, s_21_26, s_21_27, s_21_28, s_21_29, s_21_30, s_21_31, s_21_32, s_21_33, s_21_34, s_21_35, s_21_36, s_21_37, s_21_38, s_21_39, s_21_40, s_21_41, s_21_42, s_21_43, s_21_44, s_21_45, s_21_46, s_21_47, s_21_48, s_21_49, s_21_50, s_21_51, s_21_52;
    divider_cell cell_21_21(empty21, c_21_21, divisor[31], s_20_21, c_21_22, c_20_20);
    divider_cell cell_21_22(s_21_22, c_21_22, divisor[30], s_20_22, c_21_23, c_20_20);
    divider_cell cell_21_23(s_21_23, c_21_23, divisor[29], s_20_23, c_21_24, c_20_20);
    divider_cell cell_21_24(s_21_24, c_21_24, divisor[28], s_20_24, c_21_25, c_20_20);
    divider_cell cell_21_25(s_21_25, c_21_25, divisor[27], s_20_25, c_21_26, c_20_20);
    divider_cell cell_21_26(s_21_26, c_21_26, divisor[26], s_20_26, c_21_27, c_20_20);
    divider_cell cell_21_27(s_21_27, c_21_27, divisor[25], s_20_27, c_21_28, c_20_20);
    divider_cell cell_21_28(s_21_28, c_21_28, divisor[24], s_20_28, c_21_29, c_20_20);
    divider_cell cell_21_29(s_21_29, c_21_29, divisor[23], s_20_29, c_21_30, c_20_20);
    divider_cell cell_21_30(s_21_30, c_21_30, divisor[22], s_20_30, c_21_31, c_20_20);
    divider_cell cell_21_31(s_21_31, c_21_31, divisor[21], s_20_31, c_21_32, c_20_20);
    divider_cell cell_21_32(s_21_32, c_21_32, divisor[20], s_20_32, c_21_33, c_20_20);
    divider_cell cell_21_33(s_21_33, c_21_33, divisor[19], s_20_33, c_21_34, c_20_20);
    divider_cell cell_21_34(s_21_34, c_21_34, divisor[18], s_20_34, c_21_35, c_20_20);
    divider_cell cell_21_35(s_21_35, c_21_35, divisor[17], s_20_35, c_21_36, c_20_20);
    divider_cell cell_21_36(s_21_36, c_21_36, divisor[16], s_20_36, c_21_37, c_20_20);
    divider_cell cell_21_37(s_21_37, c_21_37, divisor[15], s_20_37, c_21_38, c_20_20);
    divider_cell cell_21_38(s_21_38, c_21_38, divisor[14], s_20_38, c_21_39, c_20_20);
    divider_cell cell_21_39(s_21_39, c_21_39, divisor[13], s_20_39, c_21_40, c_20_20);
    divider_cell cell_21_40(s_21_40, c_21_40, divisor[12], s_20_40, c_21_41, c_20_20);
    divider_cell cell_21_41(s_21_41, c_21_41, divisor[11], s_20_41, c_21_42, c_20_20);
    divider_cell cell_21_42(s_21_42, c_21_42, divisor[10], s_20_42, c_21_43, c_20_20);
    divider_cell cell_21_43(s_21_43, c_21_43, divisor[9], s_20_43, c_21_44, c_20_20);
    divider_cell cell_21_44(s_21_44, c_21_44, divisor[8], s_20_44, c_21_45, c_20_20);
    divider_cell cell_21_45(s_21_45, c_21_45, divisor[7], s_20_45, c_21_46, c_20_20);
    divider_cell cell_21_46(s_21_46, c_21_46, divisor[6], s_20_46, c_21_47, c_20_20);
    divider_cell cell_21_47(s_21_47, c_21_47, divisor[5], s_20_47, c_21_48, c_20_20);
    divider_cell cell_21_48(s_21_48, c_21_48, divisor[4], s_20_48, c_21_49, c_20_20);
    divider_cell cell_21_49(s_21_49, c_21_49, divisor[3], s_20_49, c_21_50, c_20_20);
    divider_cell cell_21_50(s_21_50, c_21_50, divisor[2], s_20_50, c_21_51, c_20_20);
    divider_cell cell_21_51(s_21_51, c_21_51, divisor[1], s_20_51, c_21_52, c_20_20);
    divider_cell cell_21_52(s_21_52, c_21_52, divisor[0], dividend[10], c_20_20, c_20_20);
    assign div_result[10] = c_21_21;
    wire c_22_22, c_22_23, c_22_24, c_22_25, c_22_26, c_22_27, c_22_28, c_22_29, c_22_30, c_22_31, c_22_32, c_22_33, c_22_34, c_22_35, c_22_36, c_22_37, c_22_38, c_22_39, c_22_40, c_22_41, c_22_42, c_22_43, c_22_44, c_22_45, c_22_46, c_22_47, c_22_48, c_22_49, c_22_50, c_22_51, c_22_52, c_22_53;
    wire empty22, s_22_23, s_22_24, s_22_25, s_22_26, s_22_27, s_22_28, s_22_29, s_22_30, s_22_31, s_22_32, s_22_33, s_22_34, s_22_35, s_22_36, s_22_37, s_22_38, s_22_39, s_22_40, s_22_41, s_22_42, s_22_43, s_22_44, s_22_45, s_22_46, s_22_47, s_22_48, s_22_49, s_22_50, s_22_51, s_22_52, s_22_53;
    divider_cell cell_22_22(empty22, c_22_22, divisor[31], s_21_22, c_22_23, c_21_21);
    divider_cell cell_22_23(s_22_23, c_22_23, divisor[30], s_21_23, c_22_24, c_21_21);
    divider_cell cell_22_24(s_22_24, c_22_24, divisor[29], s_21_24, c_22_25, c_21_21);
    divider_cell cell_22_25(s_22_25, c_22_25, divisor[28], s_21_25, c_22_26, c_21_21);
    divider_cell cell_22_26(s_22_26, c_22_26, divisor[27], s_21_26, c_22_27, c_21_21);
    divider_cell cell_22_27(s_22_27, c_22_27, divisor[26], s_21_27, c_22_28, c_21_21);
    divider_cell cell_22_28(s_22_28, c_22_28, divisor[25], s_21_28, c_22_29, c_21_21);
    divider_cell cell_22_29(s_22_29, c_22_29, divisor[24], s_21_29, c_22_30, c_21_21);
    divider_cell cell_22_30(s_22_30, c_22_30, divisor[23], s_21_30, c_22_31, c_21_21);
    divider_cell cell_22_31(s_22_31, c_22_31, divisor[22], s_21_31, c_22_32, c_21_21);
    divider_cell cell_22_32(s_22_32, c_22_32, divisor[21], s_21_32, c_22_33, c_21_21);
    divider_cell cell_22_33(s_22_33, c_22_33, divisor[20], s_21_33, c_22_34, c_21_21);
    divider_cell cell_22_34(s_22_34, c_22_34, divisor[19], s_21_34, c_22_35, c_21_21);
    divider_cell cell_22_35(s_22_35, c_22_35, divisor[18], s_21_35, c_22_36, c_21_21);
    divider_cell cell_22_36(s_22_36, c_22_36, divisor[17], s_21_36, c_22_37, c_21_21);
    divider_cell cell_22_37(s_22_37, c_22_37, divisor[16], s_21_37, c_22_38, c_21_21);
    divider_cell cell_22_38(s_22_38, c_22_38, divisor[15], s_21_38, c_22_39, c_21_21);
    divider_cell cell_22_39(s_22_39, c_22_39, divisor[14], s_21_39, c_22_40, c_21_21);
    divider_cell cell_22_40(s_22_40, c_22_40, divisor[13], s_21_40, c_22_41, c_21_21);
    divider_cell cell_22_41(s_22_41, c_22_41, divisor[12], s_21_41, c_22_42, c_21_21);
    divider_cell cell_22_42(s_22_42, c_22_42, divisor[11], s_21_42, c_22_43, c_21_21);
    divider_cell cell_22_43(s_22_43, c_22_43, divisor[10], s_21_43, c_22_44, c_21_21);
    divider_cell cell_22_44(s_22_44, c_22_44, divisor[9], s_21_44, c_22_45, c_21_21);
    divider_cell cell_22_45(s_22_45, c_22_45, divisor[8], s_21_45, c_22_46, c_21_21);
    divider_cell cell_22_46(s_22_46, c_22_46, divisor[7], s_21_46, c_22_47, c_21_21);
    divider_cell cell_22_47(s_22_47, c_22_47, divisor[6], s_21_47, c_22_48, c_21_21);
    divider_cell cell_22_48(s_22_48, c_22_48, divisor[5], s_21_48, c_22_49, c_21_21);
    divider_cell cell_22_49(s_22_49, c_22_49, divisor[4], s_21_49, c_22_50, c_21_21);
    divider_cell cell_22_50(s_22_50, c_22_50, divisor[3], s_21_50, c_22_51, c_21_21);
    divider_cell cell_22_51(s_22_51, c_22_51, divisor[2], s_21_51, c_22_52, c_21_21);
    divider_cell cell_22_52(s_22_52, c_22_52, divisor[1], s_21_52, c_22_53, c_21_21);
    divider_cell cell_22_53(s_22_53, c_22_53, divisor[0], dividend[9], c_21_21, c_21_21);
    assign div_result[9] = c_22_22;
    wire c_23_23, c_23_24, c_23_25, c_23_26, c_23_27, c_23_28, c_23_29, c_23_30, c_23_31, c_23_32, c_23_33, c_23_34, c_23_35, c_23_36, c_23_37, c_23_38, c_23_39, c_23_40, c_23_41, c_23_42, c_23_43, c_23_44, c_23_45, c_23_46, c_23_47, c_23_48, c_23_49, c_23_50, c_23_51, c_23_52, c_23_53, c_23_54;
    wire empty23, s_23_24, s_23_25, s_23_26, s_23_27, s_23_28, s_23_29, s_23_30, s_23_31, s_23_32, s_23_33, s_23_34, s_23_35, s_23_36, s_23_37, s_23_38, s_23_39, s_23_40, s_23_41, s_23_42, s_23_43, s_23_44, s_23_45, s_23_46, s_23_47, s_23_48, s_23_49, s_23_50, s_23_51, s_23_52, s_23_53, s_23_54;
    divider_cell cell_23_23(empty23, c_23_23, divisor[31], s_22_23, c_23_24, c_22_22);
    divider_cell cell_23_24(s_23_24, c_23_24, divisor[30], s_22_24, c_23_25, c_22_22);
    divider_cell cell_23_25(s_23_25, c_23_25, divisor[29], s_22_25, c_23_26, c_22_22);
    divider_cell cell_23_26(s_23_26, c_23_26, divisor[28], s_22_26, c_23_27, c_22_22);
    divider_cell cell_23_27(s_23_27, c_23_27, divisor[27], s_22_27, c_23_28, c_22_22);
    divider_cell cell_23_28(s_23_28, c_23_28, divisor[26], s_22_28, c_23_29, c_22_22);
    divider_cell cell_23_29(s_23_29, c_23_29, divisor[25], s_22_29, c_23_30, c_22_22);
    divider_cell cell_23_30(s_23_30, c_23_30, divisor[24], s_22_30, c_23_31, c_22_22);
    divider_cell cell_23_31(s_23_31, c_23_31, divisor[23], s_22_31, c_23_32, c_22_22);
    divider_cell cell_23_32(s_23_32, c_23_32, divisor[22], s_22_32, c_23_33, c_22_22);
    divider_cell cell_23_33(s_23_33, c_23_33, divisor[21], s_22_33, c_23_34, c_22_22);
    divider_cell cell_23_34(s_23_34, c_23_34, divisor[20], s_22_34, c_23_35, c_22_22);
    divider_cell cell_23_35(s_23_35, c_23_35, divisor[19], s_22_35, c_23_36, c_22_22);
    divider_cell cell_23_36(s_23_36, c_23_36, divisor[18], s_22_36, c_23_37, c_22_22);
    divider_cell cell_23_37(s_23_37, c_23_37, divisor[17], s_22_37, c_23_38, c_22_22);
    divider_cell cell_23_38(s_23_38, c_23_38, divisor[16], s_22_38, c_23_39, c_22_22);
    divider_cell cell_23_39(s_23_39, c_23_39, divisor[15], s_22_39, c_23_40, c_22_22);
    divider_cell cell_23_40(s_23_40, c_23_40, divisor[14], s_22_40, c_23_41, c_22_22);
    divider_cell cell_23_41(s_23_41, c_23_41, divisor[13], s_22_41, c_23_42, c_22_22);
    divider_cell cell_23_42(s_23_42, c_23_42, divisor[12], s_22_42, c_23_43, c_22_22);
    divider_cell cell_23_43(s_23_43, c_23_43, divisor[11], s_22_43, c_23_44, c_22_22);
    divider_cell cell_23_44(s_23_44, c_23_44, divisor[10], s_22_44, c_23_45, c_22_22);
    divider_cell cell_23_45(s_23_45, c_23_45, divisor[9], s_22_45, c_23_46, c_22_22);
    divider_cell cell_23_46(s_23_46, c_23_46, divisor[8], s_22_46, c_23_47, c_22_22);
    divider_cell cell_23_47(s_23_47, c_23_47, divisor[7], s_22_47, c_23_48, c_22_22);
    divider_cell cell_23_48(s_23_48, c_23_48, divisor[6], s_22_48, c_23_49, c_22_22);
    divider_cell cell_23_49(s_23_49, c_23_49, divisor[5], s_22_49, c_23_50, c_22_22);
    divider_cell cell_23_50(s_23_50, c_23_50, divisor[4], s_22_50, c_23_51, c_22_22);
    divider_cell cell_23_51(s_23_51, c_23_51, divisor[3], s_22_51, c_23_52, c_22_22);
    divider_cell cell_23_52(s_23_52, c_23_52, divisor[2], s_22_52, c_23_53, c_22_22);
    divider_cell cell_23_53(s_23_53, c_23_53, divisor[1], s_22_53, c_23_54, c_22_22);
    divider_cell cell_23_54(s_23_54, c_23_54, divisor[0], dividend[8], c_22_22, c_22_22);
    assign div_result[8] = c_23_23;
    wire c_24_24, c_24_25, c_24_26, c_24_27, c_24_28, c_24_29, c_24_30, c_24_31, c_24_32, c_24_33, c_24_34, c_24_35, c_24_36, c_24_37, c_24_38, c_24_39, c_24_40, c_24_41, c_24_42, c_24_43, c_24_44, c_24_45, c_24_46, c_24_47, c_24_48, c_24_49, c_24_50, c_24_51, c_24_52, c_24_53, c_24_54, c_24_55;
    wire empty24, s_24_25, s_24_26, s_24_27, s_24_28, s_24_29, s_24_30, s_24_31, s_24_32, s_24_33, s_24_34, s_24_35, s_24_36, s_24_37, s_24_38, s_24_39, s_24_40, s_24_41, s_24_42, s_24_43, s_24_44, s_24_45, s_24_46, s_24_47, s_24_48, s_24_49, s_24_50, s_24_51, s_24_52, s_24_53, s_24_54, s_24_55;
    divider_cell cell_24_24(empty24, c_24_24, divisor[31], s_23_24, c_24_25, c_23_23);
    divider_cell cell_24_25(s_24_25, c_24_25, divisor[30], s_23_25, c_24_26, c_23_23);
    divider_cell cell_24_26(s_24_26, c_24_26, divisor[29], s_23_26, c_24_27, c_23_23);
    divider_cell cell_24_27(s_24_27, c_24_27, divisor[28], s_23_27, c_24_28, c_23_23);
    divider_cell cell_24_28(s_24_28, c_24_28, divisor[27], s_23_28, c_24_29, c_23_23);
    divider_cell cell_24_29(s_24_29, c_24_29, divisor[26], s_23_29, c_24_30, c_23_23);
    divider_cell cell_24_30(s_24_30, c_24_30, divisor[25], s_23_30, c_24_31, c_23_23);
    divider_cell cell_24_31(s_24_31, c_24_31, divisor[24], s_23_31, c_24_32, c_23_23);
    divider_cell cell_24_32(s_24_32, c_24_32, divisor[23], s_23_32, c_24_33, c_23_23);
    divider_cell cell_24_33(s_24_33, c_24_33, divisor[22], s_23_33, c_24_34, c_23_23);
    divider_cell cell_24_34(s_24_34, c_24_34, divisor[21], s_23_34, c_24_35, c_23_23);
    divider_cell cell_24_35(s_24_35, c_24_35, divisor[20], s_23_35, c_24_36, c_23_23);
    divider_cell cell_24_36(s_24_36, c_24_36, divisor[19], s_23_36, c_24_37, c_23_23);
    divider_cell cell_24_37(s_24_37, c_24_37, divisor[18], s_23_37, c_24_38, c_23_23);
    divider_cell cell_24_38(s_24_38, c_24_38, divisor[17], s_23_38, c_24_39, c_23_23);
    divider_cell cell_24_39(s_24_39, c_24_39, divisor[16], s_23_39, c_24_40, c_23_23);
    divider_cell cell_24_40(s_24_40, c_24_40, divisor[15], s_23_40, c_24_41, c_23_23);
    divider_cell cell_24_41(s_24_41, c_24_41, divisor[14], s_23_41, c_24_42, c_23_23);
    divider_cell cell_24_42(s_24_42, c_24_42, divisor[13], s_23_42, c_24_43, c_23_23);
    divider_cell cell_24_43(s_24_43, c_24_43, divisor[12], s_23_43, c_24_44, c_23_23);
    divider_cell cell_24_44(s_24_44, c_24_44, divisor[11], s_23_44, c_24_45, c_23_23);
    divider_cell cell_24_45(s_24_45, c_24_45, divisor[10], s_23_45, c_24_46, c_23_23);
    divider_cell cell_24_46(s_24_46, c_24_46, divisor[9], s_23_46, c_24_47, c_23_23);
    divider_cell cell_24_47(s_24_47, c_24_47, divisor[8], s_23_47, c_24_48, c_23_23);
    divider_cell cell_24_48(s_24_48, c_24_48, divisor[7], s_23_48, c_24_49, c_23_23);
    divider_cell cell_24_49(s_24_49, c_24_49, divisor[6], s_23_49, c_24_50, c_23_23);
    divider_cell cell_24_50(s_24_50, c_24_50, divisor[5], s_23_50, c_24_51, c_23_23);
    divider_cell cell_24_51(s_24_51, c_24_51, divisor[4], s_23_51, c_24_52, c_23_23);
    divider_cell cell_24_52(s_24_52, c_24_52, divisor[3], s_23_52, c_24_53, c_23_23);
    divider_cell cell_24_53(s_24_53, c_24_53, divisor[2], s_23_53, c_24_54, c_23_23);
    divider_cell cell_24_54(s_24_54, c_24_54, divisor[1], s_23_54, c_24_55, c_23_23);
    divider_cell cell_24_55(s_24_55, c_24_55, divisor[0], dividend[7], c_23_23, c_23_23);
    assign div_result[7] = c_24_24;
    wire c_25_25, c_25_26, c_25_27, c_25_28, c_25_29, c_25_30, c_25_31, c_25_32, c_25_33, c_25_34, c_25_35, c_25_36, c_25_37, c_25_38, c_25_39, c_25_40, c_25_41, c_25_42, c_25_43, c_25_44, c_25_45, c_25_46, c_25_47, c_25_48, c_25_49, c_25_50, c_25_51, c_25_52, c_25_53, c_25_54, c_25_55, c_25_56;
    wire empty25, s_25_26, s_25_27, s_25_28, s_25_29, s_25_30, s_25_31, s_25_32, s_25_33, s_25_34, s_25_35, s_25_36, s_25_37, s_25_38, s_25_39, s_25_40, s_25_41, s_25_42, s_25_43, s_25_44, s_25_45, s_25_46, s_25_47, s_25_48, s_25_49, s_25_50, s_25_51, s_25_52, s_25_53, s_25_54, s_25_55, s_25_56;
    divider_cell cell_25_25(empty25, c_25_25, divisor[31], s_24_25, c_25_26, c_24_24);
    divider_cell cell_25_26(s_25_26, c_25_26, divisor[30], s_24_26, c_25_27, c_24_24);
    divider_cell cell_25_27(s_25_27, c_25_27, divisor[29], s_24_27, c_25_28, c_24_24);
    divider_cell cell_25_28(s_25_28, c_25_28, divisor[28], s_24_28, c_25_29, c_24_24);
    divider_cell cell_25_29(s_25_29, c_25_29, divisor[27], s_24_29, c_25_30, c_24_24);
    divider_cell cell_25_30(s_25_30, c_25_30, divisor[26], s_24_30, c_25_31, c_24_24);
    divider_cell cell_25_31(s_25_31, c_25_31, divisor[25], s_24_31, c_25_32, c_24_24);
    divider_cell cell_25_32(s_25_32, c_25_32, divisor[24], s_24_32, c_25_33, c_24_24);
    divider_cell cell_25_33(s_25_33, c_25_33, divisor[23], s_24_33, c_25_34, c_24_24);
    divider_cell cell_25_34(s_25_34, c_25_34, divisor[22], s_24_34, c_25_35, c_24_24);
    divider_cell cell_25_35(s_25_35, c_25_35, divisor[21], s_24_35, c_25_36, c_24_24);
    divider_cell cell_25_36(s_25_36, c_25_36, divisor[20], s_24_36, c_25_37, c_24_24);
    divider_cell cell_25_37(s_25_37, c_25_37, divisor[19], s_24_37, c_25_38, c_24_24);
    divider_cell cell_25_38(s_25_38, c_25_38, divisor[18], s_24_38, c_25_39, c_24_24);
    divider_cell cell_25_39(s_25_39, c_25_39, divisor[17], s_24_39, c_25_40, c_24_24);
    divider_cell cell_25_40(s_25_40, c_25_40, divisor[16], s_24_40, c_25_41, c_24_24);
    divider_cell cell_25_41(s_25_41, c_25_41, divisor[15], s_24_41, c_25_42, c_24_24);
    divider_cell cell_25_42(s_25_42, c_25_42, divisor[14], s_24_42, c_25_43, c_24_24);
    divider_cell cell_25_43(s_25_43, c_25_43, divisor[13], s_24_43, c_25_44, c_24_24);
    divider_cell cell_25_44(s_25_44, c_25_44, divisor[12], s_24_44, c_25_45, c_24_24);
    divider_cell cell_25_45(s_25_45, c_25_45, divisor[11], s_24_45, c_25_46, c_24_24);
    divider_cell cell_25_46(s_25_46, c_25_46, divisor[10], s_24_46, c_25_47, c_24_24);
    divider_cell cell_25_47(s_25_47, c_25_47, divisor[9], s_24_47, c_25_48, c_24_24);
    divider_cell cell_25_48(s_25_48, c_25_48, divisor[8], s_24_48, c_25_49, c_24_24);
    divider_cell cell_25_49(s_25_49, c_25_49, divisor[7], s_24_49, c_25_50, c_24_24);
    divider_cell cell_25_50(s_25_50, c_25_50, divisor[6], s_24_50, c_25_51, c_24_24);
    divider_cell cell_25_51(s_25_51, c_25_51, divisor[5], s_24_51, c_25_52, c_24_24);
    divider_cell cell_25_52(s_25_52, c_25_52, divisor[4], s_24_52, c_25_53, c_24_24);
    divider_cell cell_25_53(s_25_53, c_25_53, divisor[3], s_24_53, c_25_54, c_24_24);
    divider_cell cell_25_54(s_25_54, c_25_54, divisor[2], s_24_54, c_25_55, c_24_24);
    divider_cell cell_25_55(s_25_55, c_25_55, divisor[1], s_24_55, c_25_56, c_24_24);
    divider_cell cell_25_56(s_25_56, c_25_56, divisor[0], dividend[6], c_24_24, c_24_24);
    assign div_result[6] = c_25_25;
    wire c_26_26, c_26_27, c_26_28, c_26_29, c_26_30, c_26_31, c_26_32, c_26_33, c_26_34, c_26_35, c_26_36, c_26_37, c_26_38, c_26_39, c_26_40, c_26_41, c_26_42, c_26_43, c_26_44, c_26_45, c_26_46, c_26_47, c_26_48, c_26_49, c_26_50, c_26_51, c_26_52, c_26_53, c_26_54, c_26_55, c_26_56, c_26_57;
    wire empty26, s_26_27, s_26_28, s_26_29, s_26_30, s_26_31, s_26_32, s_26_33, s_26_34, s_26_35, s_26_36, s_26_37, s_26_38, s_26_39, s_26_40, s_26_41, s_26_42, s_26_43, s_26_44, s_26_45, s_26_46, s_26_47, s_26_48, s_26_49, s_26_50, s_26_51, s_26_52, s_26_53, s_26_54, s_26_55, s_26_56, s_26_57;
    divider_cell cell_26_26(empty26, c_26_26, divisor[31], s_25_26, c_26_27, c_25_25);
    divider_cell cell_26_27(s_26_27, c_26_27, divisor[30], s_25_27, c_26_28, c_25_25);
    divider_cell cell_26_28(s_26_28, c_26_28, divisor[29], s_25_28, c_26_29, c_25_25);
    divider_cell cell_26_29(s_26_29, c_26_29, divisor[28], s_25_29, c_26_30, c_25_25);
    divider_cell cell_26_30(s_26_30, c_26_30, divisor[27], s_25_30, c_26_31, c_25_25);
    divider_cell cell_26_31(s_26_31, c_26_31, divisor[26], s_25_31, c_26_32, c_25_25);
    divider_cell cell_26_32(s_26_32, c_26_32, divisor[25], s_25_32, c_26_33, c_25_25);
    divider_cell cell_26_33(s_26_33, c_26_33, divisor[24], s_25_33, c_26_34, c_25_25);
    divider_cell cell_26_34(s_26_34, c_26_34, divisor[23], s_25_34, c_26_35, c_25_25);
    divider_cell cell_26_35(s_26_35, c_26_35, divisor[22], s_25_35, c_26_36, c_25_25);
    divider_cell cell_26_36(s_26_36, c_26_36, divisor[21], s_25_36, c_26_37, c_25_25);
    divider_cell cell_26_37(s_26_37, c_26_37, divisor[20], s_25_37, c_26_38, c_25_25);
    divider_cell cell_26_38(s_26_38, c_26_38, divisor[19], s_25_38, c_26_39, c_25_25);
    divider_cell cell_26_39(s_26_39, c_26_39, divisor[18], s_25_39, c_26_40, c_25_25);
    divider_cell cell_26_40(s_26_40, c_26_40, divisor[17], s_25_40, c_26_41, c_25_25);
    divider_cell cell_26_41(s_26_41, c_26_41, divisor[16], s_25_41, c_26_42, c_25_25);
    divider_cell cell_26_42(s_26_42, c_26_42, divisor[15], s_25_42, c_26_43, c_25_25);
    divider_cell cell_26_43(s_26_43, c_26_43, divisor[14], s_25_43, c_26_44, c_25_25);
    divider_cell cell_26_44(s_26_44, c_26_44, divisor[13], s_25_44, c_26_45, c_25_25);
    divider_cell cell_26_45(s_26_45, c_26_45, divisor[12], s_25_45, c_26_46, c_25_25);
    divider_cell cell_26_46(s_26_46, c_26_46, divisor[11], s_25_46, c_26_47, c_25_25);
    divider_cell cell_26_47(s_26_47, c_26_47, divisor[10], s_25_47, c_26_48, c_25_25);
    divider_cell cell_26_48(s_26_48, c_26_48, divisor[9], s_25_48, c_26_49, c_25_25);
    divider_cell cell_26_49(s_26_49, c_26_49, divisor[8], s_25_49, c_26_50, c_25_25);
    divider_cell cell_26_50(s_26_50, c_26_50, divisor[7], s_25_50, c_26_51, c_25_25);
    divider_cell cell_26_51(s_26_51, c_26_51, divisor[6], s_25_51, c_26_52, c_25_25);
    divider_cell cell_26_52(s_26_52, c_26_52, divisor[5], s_25_52, c_26_53, c_25_25);
    divider_cell cell_26_53(s_26_53, c_26_53, divisor[4], s_25_53, c_26_54, c_25_25);
    divider_cell cell_26_54(s_26_54, c_26_54, divisor[3], s_25_54, c_26_55, c_25_25);
    divider_cell cell_26_55(s_26_55, c_26_55, divisor[2], s_25_55, c_26_56, c_25_25);
    divider_cell cell_26_56(s_26_56, c_26_56, divisor[1], s_25_56, c_26_57, c_25_25);
    divider_cell cell_26_57(s_26_57, c_26_57, divisor[0], dividend[5], c_25_25, c_25_25);
    assign div_result[5] = c_26_26;
    wire c_27_27, c_27_28, c_27_29, c_27_30, c_27_31, c_27_32, c_27_33, c_27_34, c_27_35, c_27_36, c_27_37, c_27_38, c_27_39, c_27_40, c_27_41, c_27_42, c_27_43, c_27_44, c_27_45, c_27_46, c_27_47, c_27_48, c_27_49, c_27_50, c_27_51, c_27_52, c_27_53, c_27_54, c_27_55, c_27_56, c_27_57, c_27_58;
    wire empty27, s_27_28, s_27_29, s_27_30, s_27_31, s_27_32, s_27_33, s_27_34, s_27_35, s_27_36, s_27_37, s_27_38, s_27_39, s_27_40, s_27_41, s_27_42, s_27_43, s_27_44, s_27_45, s_27_46, s_27_47, s_27_48, s_27_49, s_27_50, s_27_51, s_27_52, s_27_53, s_27_54, s_27_55, s_27_56, s_27_57, s_27_58;
    divider_cell cell_27_27(empty27, c_27_27, divisor[31], s_26_27, c_27_28, c_26_26);
    divider_cell cell_27_28(s_27_28, c_27_28, divisor[30], s_26_28, c_27_29, c_26_26);
    divider_cell cell_27_29(s_27_29, c_27_29, divisor[29], s_26_29, c_27_30, c_26_26);
    divider_cell cell_27_30(s_27_30, c_27_30, divisor[28], s_26_30, c_27_31, c_26_26);
    divider_cell cell_27_31(s_27_31, c_27_31, divisor[27], s_26_31, c_27_32, c_26_26);
    divider_cell cell_27_32(s_27_32, c_27_32, divisor[26], s_26_32, c_27_33, c_26_26);
    divider_cell cell_27_33(s_27_33, c_27_33, divisor[25], s_26_33, c_27_34, c_26_26);
    divider_cell cell_27_34(s_27_34, c_27_34, divisor[24], s_26_34, c_27_35, c_26_26);
    divider_cell cell_27_35(s_27_35, c_27_35, divisor[23], s_26_35, c_27_36, c_26_26);
    divider_cell cell_27_36(s_27_36, c_27_36, divisor[22], s_26_36, c_27_37, c_26_26);
    divider_cell cell_27_37(s_27_37, c_27_37, divisor[21], s_26_37, c_27_38, c_26_26);
    divider_cell cell_27_38(s_27_38, c_27_38, divisor[20], s_26_38, c_27_39, c_26_26);
    divider_cell cell_27_39(s_27_39, c_27_39, divisor[19], s_26_39, c_27_40, c_26_26);
    divider_cell cell_27_40(s_27_40, c_27_40, divisor[18], s_26_40, c_27_41, c_26_26);
    divider_cell cell_27_41(s_27_41, c_27_41, divisor[17], s_26_41, c_27_42, c_26_26);
    divider_cell cell_27_42(s_27_42, c_27_42, divisor[16], s_26_42, c_27_43, c_26_26);
    divider_cell cell_27_43(s_27_43, c_27_43, divisor[15], s_26_43, c_27_44, c_26_26);
    divider_cell cell_27_44(s_27_44, c_27_44, divisor[14], s_26_44, c_27_45, c_26_26);
    divider_cell cell_27_45(s_27_45, c_27_45, divisor[13], s_26_45, c_27_46, c_26_26);
    divider_cell cell_27_46(s_27_46, c_27_46, divisor[12], s_26_46, c_27_47, c_26_26);
    divider_cell cell_27_47(s_27_47, c_27_47, divisor[11], s_26_47, c_27_48, c_26_26);
    divider_cell cell_27_48(s_27_48, c_27_48, divisor[10], s_26_48, c_27_49, c_26_26);
    divider_cell cell_27_49(s_27_49, c_27_49, divisor[9], s_26_49, c_27_50, c_26_26);
    divider_cell cell_27_50(s_27_50, c_27_50, divisor[8], s_26_50, c_27_51, c_26_26);
    divider_cell cell_27_51(s_27_51, c_27_51, divisor[7], s_26_51, c_27_52, c_26_26);
    divider_cell cell_27_52(s_27_52, c_27_52, divisor[6], s_26_52, c_27_53, c_26_26);
    divider_cell cell_27_53(s_27_53, c_27_53, divisor[5], s_26_53, c_27_54, c_26_26);
    divider_cell cell_27_54(s_27_54, c_27_54, divisor[4], s_26_54, c_27_55, c_26_26);
    divider_cell cell_27_55(s_27_55, c_27_55, divisor[3], s_26_55, c_27_56, c_26_26);
    divider_cell cell_27_56(s_27_56, c_27_56, divisor[2], s_26_56, c_27_57, c_26_26);
    divider_cell cell_27_57(s_27_57, c_27_57, divisor[1], s_26_57, c_27_58, c_26_26);
    divider_cell cell_27_58(s_27_58, c_27_58, divisor[0], dividend[4], c_26_26, c_26_26);
    assign div_result[4] = c_27_27;
    wire c_28_28, c_28_29, c_28_30, c_28_31, c_28_32, c_28_33, c_28_34, c_28_35, c_28_36, c_28_37, c_28_38, c_28_39, c_28_40, c_28_41, c_28_42, c_28_43, c_28_44, c_28_45, c_28_46, c_28_47, c_28_48, c_28_49, c_28_50, c_28_51, c_28_52, c_28_53, c_28_54, c_28_55, c_28_56, c_28_57, c_28_58, c_28_59;
    wire empty28, s_28_29, s_28_30, s_28_31, s_28_32, s_28_33, s_28_34, s_28_35, s_28_36, s_28_37, s_28_38, s_28_39, s_28_40, s_28_41, s_28_42, s_28_43, s_28_44, s_28_45, s_28_46, s_28_47, s_28_48, s_28_49, s_28_50, s_28_51, s_28_52, s_28_53, s_28_54, s_28_55, s_28_56, s_28_57, s_28_58, s_28_59;
    divider_cell cell_28_28(empty28, c_28_28, divisor[31], s_27_28, c_28_29, c_27_27);
    divider_cell cell_28_29(s_28_29, c_28_29, divisor[30], s_27_29, c_28_30, c_27_27);
    divider_cell cell_28_30(s_28_30, c_28_30, divisor[29], s_27_30, c_28_31, c_27_27);
    divider_cell cell_28_31(s_28_31, c_28_31, divisor[28], s_27_31, c_28_32, c_27_27);
    divider_cell cell_28_32(s_28_32, c_28_32, divisor[27], s_27_32, c_28_33, c_27_27);
    divider_cell cell_28_33(s_28_33, c_28_33, divisor[26], s_27_33, c_28_34, c_27_27);
    divider_cell cell_28_34(s_28_34, c_28_34, divisor[25], s_27_34, c_28_35, c_27_27);
    divider_cell cell_28_35(s_28_35, c_28_35, divisor[24], s_27_35, c_28_36, c_27_27);
    divider_cell cell_28_36(s_28_36, c_28_36, divisor[23], s_27_36, c_28_37, c_27_27);
    divider_cell cell_28_37(s_28_37, c_28_37, divisor[22], s_27_37, c_28_38, c_27_27);
    divider_cell cell_28_38(s_28_38, c_28_38, divisor[21], s_27_38, c_28_39, c_27_27);
    divider_cell cell_28_39(s_28_39, c_28_39, divisor[20], s_27_39, c_28_40, c_27_27);
    divider_cell cell_28_40(s_28_40, c_28_40, divisor[19], s_27_40, c_28_41, c_27_27);
    divider_cell cell_28_41(s_28_41, c_28_41, divisor[18], s_27_41, c_28_42, c_27_27);
    divider_cell cell_28_42(s_28_42, c_28_42, divisor[17], s_27_42, c_28_43, c_27_27);
    divider_cell cell_28_43(s_28_43, c_28_43, divisor[16], s_27_43, c_28_44, c_27_27);
    divider_cell cell_28_44(s_28_44, c_28_44, divisor[15], s_27_44, c_28_45, c_27_27);
    divider_cell cell_28_45(s_28_45, c_28_45, divisor[14], s_27_45, c_28_46, c_27_27);
    divider_cell cell_28_46(s_28_46, c_28_46, divisor[13], s_27_46, c_28_47, c_27_27);
    divider_cell cell_28_47(s_28_47, c_28_47, divisor[12], s_27_47, c_28_48, c_27_27);
    divider_cell cell_28_48(s_28_48, c_28_48, divisor[11], s_27_48, c_28_49, c_27_27);
    divider_cell cell_28_49(s_28_49, c_28_49, divisor[10], s_27_49, c_28_50, c_27_27);
    divider_cell cell_28_50(s_28_50, c_28_50, divisor[9], s_27_50, c_28_51, c_27_27);
    divider_cell cell_28_51(s_28_51, c_28_51, divisor[8], s_27_51, c_28_52, c_27_27);
    divider_cell cell_28_52(s_28_52, c_28_52, divisor[7], s_27_52, c_28_53, c_27_27);
    divider_cell cell_28_53(s_28_53, c_28_53, divisor[6], s_27_53, c_28_54, c_27_27);
    divider_cell cell_28_54(s_28_54, c_28_54, divisor[5], s_27_54, c_28_55, c_27_27);
    divider_cell cell_28_55(s_28_55, c_28_55, divisor[4], s_27_55, c_28_56, c_27_27);
    divider_cell cell_28_56(s_28_56, c_28_56, divisor[3], s_27_56, c_28_57, c_27_27);
    divider_cell cell_28_57(s_28_57, c_28_57, divisor[2], s_27_57, c_28_58, c_27_27);
    divider_cell cell_28_58(s_28_58, c_28_58, divisor[1], s_27_58, c_28_59, c_27_27);
    divider_cell cell_28_59(s_28_59, c_28_59, divisor[0], dividend[3], c_27_27, c_27_27);
    assign div_result[3] = c_28_28;
    wire c_29_29, c_29_30, c_29_31, c_29_32, c_29_33, c_29_34, c_29_35, c_29_36, c_29_37, c_29_38, c_29_39, c_29_40, c_29_41, c_29_42, c_29_43, c_29_44, c_29_45, c_29_46, c_29_47, c_29_48, c_29_49, c_29_50, c_29_51, c_29_52, c_29_53, c_29_54, c_29_55, c_29_56, c_29_57, c_29_58, c_29_59, c_29_60;
    wire empty29, s_29_30, s_29_31, s_29_32, s_29_33, s_29_34, s_29_35, s_29_36, s_29_37, s_29_38, s_29_39, s_29_40, s_29_41, s_29_42, s_29_43, s_29_44, s_29_45, s_29_46, s_29_47, s_29_48, s_29_49, s_29_50, s_29_51, s_29_52, s_29_53, s_29_54, s_29_55, s_29_56, s_29_57, s_29_58, s_29_59, s_29_60;
    divider_cell cell_29_29(empty29, c_29_29, divisor[31], s_28_29, c_29_30, c_28_28);
    divider_cell cell_29_30(s_29_30, c_29_30, divisor[30], s_28_30, c_29_31, c_28_28);
    divider_cell cell_29_31(s_29_31, c_29_31, divisor[29], s_28_31, c_29_32, c_28_28);
    divider_cell cell_29_32(s_29_32, c_29_32, divisor[28], s_28_32, c_29_33, c_28_28);
    divider_cell cell_29_33(s_29_33, c_29_33, divisor[27], s_28_33, c_29_34, c_28_28);
    divider_cell cell_29_34(s_29_34, c_29_34, divisor[26], s_28_34, c_29_35, c_28_28);
    divider_cell cell_29_35(s_29_35, c_29_35, divisor[25], s_28_35, c_29_36, c_28_28);
    divider_cell cell_29_36(s_29_36, c_29_36, divisor[24], s_28_36, c_29_37, c_28_28);
    divider_cell cell_29_37(s_29_37, c_29_37, divisor[23], s_28_37, c_29_38, c_28_28);
    divider_cell cell_29_38(s_29_38, c_29_38, divisor[22], s_28_38, c_29_39, c_28_28);
    divider_cell cell_29_39(s_29_39, c_29_39, divisor[21], s_28_39, c_29_40, c_28_28);
    divider_cell cell_29_40(s_29_40, c_29_40, divisor[20], s_28_40, c_29_41, c_28_28);
    divider_cell cell_29_41(s_29_41, c_29_41, divisor[19], s_28_41, c_29_42, c_28_28);
    divider_cell cell_29_42(s_29_42, c_29_42, divisor[18], s_28_42, c_29_43, c_28_28);
    divider_cell cell_29_43(s_29_43, c_29_43, divisor[17], s_28_43, c_29_44, c_28_28);
    divider_cell cell_29_44(s_29_44, c_29_44, divisor[16], s_28_44, c_29_45, c_28_28);
    divider_cell cell_29_45(s_29_45, c_29_45, divisor[15], s_28_45, c_29_46, c_28_28);
    divider_cell cell_29_46(s_29_46, c_29_46, divisor[14], s_28_46, c_29_47, c_28_28);
    divider_cell cell_29_47(s_29_47, c_29_47, divisor[13], s_28_47, c_29_48, c_28_28);
    divider_cell cell_29_48(s_29_48, c_29_48, divisor[12], s_28_48, c_29_49, c_28_28);
    divider_cell cell_29_49(s_29_49, c_29_49, divisor[11], s_28_49, c_29_50, c_28_28);
    divider_cell cell_29_50(s_29_50, c_29_50, divisor[10], s_28_50, c_29_51, c_28_28);
    divider_cell cell_29_51(s_29_51, c_29_51, divisor[9], s_28_51, c_29_52, c_28_28);
    divider_cell cell_29_52(s_29_52, c_29_52, divisor[8], s_28_52, c_29_53, c_28_28);
    divider_cell cell_29_53(s_29_53, c_29_53, divisor[7], s_28_53, c_29_54, c_28_28);
    divider_cell cell_29_54(s_29_54, c_29_54, divisor[6], s_28_54, c_29_55, c_28_28);
    divider_cell cell_29_55(s_29_55, c_29_55, divisor[5], s_28_55, c_29_56, c_28_28);
    divider_cell cell_29_56(s_29_56, c_29_56, divisor[4], s_28_56, c_29_57, c_28_28);
    divider_cell cell_29_57(s_29_57, c_29_57, divisor[3], s_28_57, c_29_58, c_28_28);
    divider_cell cell_29_58(s_29_58, c_29_58, divisor[2], s_28_58, c_29_59, c_28_28);
    divider_cell cell_29_59(s_29_59, c_29_59, divisor[1], s_28_59, c_29_60, c_28_28);
    divider_cell cell_29_60(s_29_60, c_29_60, divisor[0], dividend[2], c_28_28, c_28_28);
    assign div_result[2] = c_29_29;
    wire c_30_30, c_30_31, c_30_32, c_30_33, c_30_34, c_30_35, c_30_36, c_30_37, c_30_38, c_30_39, c_30_40, c_30_41, c_30_42, c_30_43, c_30_44, c_30_45, c_30_46, c_30_47, c_30_48, c_30_49, c_30_50, c_30_51, c_30_52, c_30_53, c_30_54, c_30_55, c_30_56, c_30_57, c_30_58, c_30_59, c_30_60, c_30_61;
    wire empty30, s_30_31, s_30_32, s_30_33, s_30_34, s_30_35, s_30_36, s_30_37, s_30_38, s_30_39, s_30_40, s_30_41, s_30_42, s_30_43, s_30_44, s_30_45, s_30_46, s_30_47, s_30_48, s_30_49, s_30_50, s_30_51, s_30_52, s_30_53, s_30_54, s_30_55, s_30_56, s_30_57, s_30_58, s_30_59, s_30_60, s_30_61;
    divider_cell cell_30_30(empty30, c_30_30, divisor[31], s_29_30, c_30_31, c_29_29);
    divider_cell cell_30_31(s_30_31, c_30_31, divisor[30], s_29_31, c_30_32, c_29_29);
    divider_cell cell_30_32(s_30_32, c_30_32, divisor[29], s_29_32, c_30_33, c_29_29);
    divider_cell cell_30_33(s_30_33, c_30_33, divisor[28], s_29_33, c_30_34, c_29_29);
    divider_cell cell_30_34(s_30_34, c_30_34, divisor[27], s_29_34, c_30_35, c_29_29);
    divider_cell cell_30_35(s_30_35, c_30_35, divisor[26], s_29_35, c_30_36, c_29_29);
    divider_cell cell_30_36(s_30_36, c_30_36, divisor[25], s_29_36, c_30_37, c_29_29);
    divider_cell cell_30_37(s_30_37, c_30_37, divisor[24], s_29_37, c_30_38, c_29_29);
    divider_cell cell_30_38(s_30_38, c_30_38, divisor[23], s_29_38, c_30_39, c_29_29);
    divider_cell cell_30_39(s_30_39, c_30_39, divisor[22], s_29_39, c_30_40, c_29_29);
    divider_cell cell_30_40(s_30_40, c_30_40, divisor[21], s_29_40, c_30_41, c_29_29);
    divider_cell cell_30_41(s_30_41, c_30_41, divisor[20], s_29_41, c_30_42, c_29_29);
    divider_cell cell_30_42(s_30_42, c_30_42, divisor[19], s_29_42, c_30_43, c_29_29);
    divider_cell cell_30_43(s_30_43, c_30_43, divisor[18], s_29_43, c_30_44, c_29_29);
    divider_cell cell_30_44(s_30_44, c_30_44, divisor[17], s_29_44, c_30_45, c_29_29);
    divider_cell cell_30_45(s_30_45, c_30_45, divisor[16], s_29_45, c_30_46, c_29_29);
    divider_cell cell_30_46(s_30_46, c_30_46, divisor[15], s_29_46, c_30_47, c_29_29);
    divider_cell cell_30_47(s_30_47, c_30_47, divisor[14], s_29_47, c_30_48, c_29_29);
    divider_cell cell_30_48(s_30_48, c_30_48, divisor[13], s_29_48, c_30_49, c_29_29);
    divider_cell cell_30_49(s_30_49, c_30_49, divisor[12], s_29_49, c_30_50, c_29_29);
    divider_cell cell_30_50(s_30_50, c_30_50, divisor[11], s_29_50, c_30_51, c_29_29);
    divider_cell cell_30_51(s_30_51, c_30_51, divisor[10], s_29_51, c_30_52, c_29_29);
    divider_cell cell_30_52(s_30_52, c_30_52, divisor[9], s_29_52, c_30_53, c_29_29);
    divider_cell cell_30_53(s_30_53, c_30_53, divisor[8], s_29_53, c_30_54, c_29_29);
    divider_cell cell_30_54(s_30_54, c_30_54, divisor[7], s_29_54, c_30_55, c_29_29);
    divider_cell cell_30_55(s_30_55, c_30_55, divisor[6], s_29_55, c_30_56, c_29_29);
    divider_cell cell_30_56(s_30_56, c_30_56, divisor[5], s_29_56, c_30_57, c_29_29);
    divider_cell cell_30_57(s_30_57, c_30_57, divisor[4], s_29_57, c_30_58, c_29_29);
    divider_cell cell_30_58(s_30_58, c_30_58, divisor[3], s_29_58, c_30_59, c_29_29);
    divider_cell cell_30_59(s_30_59, c_30_59, divisor[2], s_29_59, c_30_60, c_29_29);
    divider_cell cell_30_60(s_30_60, c_30_60, divisor[1], s_29_60, c_30_61, c_29_29);
    divider_cell cell_30_61(s_30_61, c_30_61, divisor[0], dividend[1], c_29_29, c_29_29);
    assign div_result[1] = c_30_30;
    wire c_31_31, c_31_32, c_31_33, c_31_34, c_31_35, c_31_36, c_31_37, c_31_38, c_31_39, c_31_40, c_31_41, c_31_42, c_31_43, c_31_44, c_31_45, c_31_46, c_31_47, c_31_48, c_31_49, c_31_50, c_31_51, c_31_52, c_31_53, c_31_54, c_31_55, c_31_56, c_31_57, c_31_58, c_31_59, c_31_60, c_31_61, c_31_62;
    wire empty31, s_31_32, s_31_33, s_31_34, s_31_35, s_31_36, s_31_37, s_31_38, s_31_39, s_31_40, s_31_41, s_31_42, s_31_43, s_31_44, s_31_45, s_31_46, s_31_47, s_31_48, s_31_49, s_31_50, s_31_51, s_31_52, s_31_53, s_31_54, s_31_55, s_31_56, s_31_57, s_31_58, s_31_59, s_31_60, s_31_61, s_31_62;
    divider_cell cell_31_31(empty31, c_31_31, divisor[31], s_30_31, c_31_32, c_30_30);
    divider_cell cell_31_32(s_31_32, c_31_32, divisor[30], s_30_32, c_31_33, c_30_30);
    divider_cell cell_31_33(s_31_33, c_31_33, divisor[29], s_30_33, c_31_34, c_30_30);
    divider_cell cell_31_34(s_31_34, c_31_34, divisor[28], s_30_34, c_31_35, c_30_30);
    divider_cell cell_31_35(s_31_35, c_31_35, divisor[27], s_30_35, c_31_36, c_30_30);
    divider_cell cell_31_36(s_31_36, c_31_36, divisor[26], s_30_36, c_31_37, c_30_30);
    divider_cell cell_31_37(s_31_37, c_31_37, divisor[25], s_30_37, c_31_38, c_30_30);
    divider_cell cell_31_38(s_31_38, c_31_38, divisor[24], s_30_38, c_31_39, c_30_30);
    divider_cell cell_31_39(s_31_39, c_31_39, divisor[23], s_30_39, c_31_40, c_30_30);
    divider_cell cell_31_40(s_31_40, c_31_40, divisor[22], s_30_40, c_31_41, c_30_30);
    divider_cell cell_31_41(s_31_41, c_31_41, divisor[21], s_30_41, c_31_42, c_30_30);
    divider_cell cell_31_42(s_31_42, c_31_42, divisor[20], s_30_42, c_31_43, c_30_30);
    divider_cell cell_31_43(s_31_43, c_31_43, divisor[19], s_30_43, c_31_44, c_30_30);
    divider_cell cell_31_44(s_31_44, c_31_44, divisor[18], s_30_44, c_31_45, c_30_30);
    divider_cell cell_31_45(s_31_45, c_31_45, divisor[17], s_30_45, c_31_46, c_30_30);
    divider_cell cell_31_46(s_31_46, c_31_46, divisor[16], s_30_46, c_31_47, c_30_30);
    divider_cell cell_31_47(s_31_47, c_31_47, divisor[15], s_30_47, c_31_48, c_30_30);
    divider_cell cell_31_48(s_31_48, c_31_48, divisor[14], s_30_48, c_31_49, c_30_30);
    divider_cell cell_31_49(s_31_49, c_31_49, divisor[13], s_30_49, c_31_50, c_30_30);
    divider_cell cell_31_50(s_31_50, c_31_50, divisor[12], s_30_50, c_31_51, c_30_30);
    divider_cell cell_31_51(s_31_51, c_31_51, divisor[11], s_30_51, c_31_52, c_30_30);
    divider_cell cell_31_52(s_31_52, c_31_52, divisor[10], s_30_52, c_31_53, c_30_30);
    divider_cell cell_31_53(s_31_53, c_31_53, divisor[9], s_30_53, c_31_54, c_30_30);
    divider_cell cell_31_54(s_31_54, c_31_54, divisor[8], s_30_54, c_31_55, c_30_30);
    divider_cell cell_31_55(s_31_55, c_31_55, divisor[7], s_30_55, c_31_56, c_30_30);
    divider_cell cell_31_56(s_31_56, c_31_56, divisor[6], s_30_56, c_31_57, c_30_30);
    divider_cell cell_31_57(s_31_57, c_31_57, divisor[5], s_30_57, c_31_58, c_30_30);
    divider_cell cell_31_58(s_31_58, c_31_58, divisor[4], s_30_58, c_31_59, c_30_30);
    divider_cell cell_31_59(s_31_59, c_31_59, divisor[3], s_30_59, c_31_60, c_30_30);
    divider_cell cell_31_60(s_31_60, c_31_60, divisor[2], s_30_60, c_31_61, c_30_30);
    divider_cell cell_31_61(s_31_61, c_31_61, divisor[1], s_30_61, c_31_62, c_30_30);
    divider_cell cell_31_62(s_31_62, c_31_62, divisor[0], dividend[0], c_30_30, c_30_30);
    assign div_result[0] = c_31_31;





endmodule