`timescale 1ns / 1ps
module RAM #( parameter DATA_WIDTH = 32, ADDRESS_WIDTH = 15, DEPTH = 32768) ( // //12 4096, 18 262144
    input wire                     clk,                     
    input wire                     wEn,
    // input wire                     big,
    input wire [ADDRESS_WIDTH-1:0] addr,
    input wire [DATA_WIDTH-1:0]    dataIn,
    output reg [DATA_WIDTH-1:0]    dataOut = 0);
    
    reg[DATA_WIDTH-1:0] MemoryArray[0:DEPTH-1];
    
    integer i;
    initial begin
        for (i = 0; i < DEPTH; i = i + 1) begin
            MemoryArray[i] <= 0;
        end
        // if(MEMFILE > 0) begin
        //     $readmemh(MEMFILE, MemoryArray);
        // end
    end
    
    always @(posedge clk) begin
        if(wEn) begin
            MemoryArray[addr] <= dataIn;
        end else begin
            dataOut <= MemoryArray[addr];
        end
    end

    // integer j;
    // always @(posedge (clk && big)) begin
    //     if(wEn) begin
    //         for (j = 0; j< BRAIN_SIZE; j = j+1) begin
    //             MemoryArray[addr+j] <= MemoryArray[dataIn+j]; //for loop to copy brains over very quickly
    //         end
    //     end
    // end


endmodule
