module wallace_tree_32b(result, data_operandA, data_operandB);

    input [31:0] data_operandA, data_operandB;
    output [63:0] result;

    wire w_0_0, w_0_1, w_0_2, w_0_3, w_0_4, w_0_5, w_0_6, w_0_7, w_0_8, w_0_9, w_0_10, w_0_11, w_0_12, w_0_13, w_0_14, w_0_15, w_0_16, w_0_17, w_0_18, w_0_19, w_0_20, w_0_21, w_0_22, w_0_23, w_0_24, w_0_25, w_0_26, w_0_27, w_0_28, w_0_29, w_0_30, w_0_31;
    assign w_0_0 = data_operandA[0] & data_operandB[0];
    assign w_0_1 = data_operandA[1] & data_operandB[0];
    assign w_0_2 = data_operandA[2] & data_operandB[0];
    assign w_0_3 = data_operandA[3] & data_operandB[0];
    assign w_0_4 = data_operandA[4] & data_operandB[0];
    assign w_0_5 = data_operandA[5] & data_operandB[0];
    assign w_0_6 = data_operandA[6] & data_operandB[0];
    assign w_0_7 = data_operandA[7] & data_operandB[0];
    assign w_0_8 = data_operandA[8] & data_operandB[0];
    assign w_0_9 = data_operandA[9] & data_operandB[0];
    assign w_0_10 = data_operandA[10] & data_operandB[0];
    assign w_0_11 = data_operandA[11] & data_operandB[0];
    assign w_0_12 = data_operandA[12] & data_operandB[0];
    assign w_0_13 = data_operandA[13] & data_operandB[0];
    assign w_0_14 = data_operandA[14] & data_operandB[0];
    assign w_0_15 = data_operandA[15] & data_operandB[0];
    assign w_0_16 = data_operandA[16] & data_operandB[0];
    assign w_0_17 = data_operandA[17] & data_operandB[0];
    assign w_0_18 = data_operandA[18] & data_operandB[0];
    assign w_0_19 = data_operandA[19] & data_operandB[0];
    assign w_0_20 = data_operandA[20] & data_operandB[0];
    assign w_0_21 = data_operandA[21] & data_operandB[0];
    assign w_0_22 = data_operandA[22] & data_operandB[0];
    assign w_0_23 = data_operandA[23] & data_operandB[0];
    assign w_0_24 = data_operandA[24] & data_operandB[0];
    assign w_0_25 = data_operandA[25] & data_operandB[0];
    assign w_0_26 = data_operandA[26] & data_operandB[0];
    assign w_0_27 = data_operandA[27] & data_operandB[0];
    assign w_0_28 = data_operandA[28] & data_operandB[0];
    assign w_0_29 = data_operandA[29] & data_operandB[0];
    assign w_0_30 = data_operandA[30] & data_operandB[0];
    assign w_0_31 = ~(data_operandA[31] & data_operandB[0]);
    assign result[0] = w_0_0;
    wire w_1_1, w_1_2, w_1_3, w_1_4, w_1_5, w_1_6, w_1_7, w_1_8, w_1_9, w_1_10, w_1_11, w_1_12, w_1_13, w_1_14, w_1_15, w_1_16, w_1_17, w_1_18, w_1_19, w_1_20, w_1_21, w_1_22, w_1_23, w_1_24, w_1_25, w_1_26, w_1_27, w_1_28, w_1_29, w_1_30, w_1_31, w_1_32;
    wire s_1_1, s_1_2, s_1_3, s_1_4, s_1_5, s_1_6, s_1_7, s_1_8, s_1_9, s_1_10, s_1_11, s_1_12, s_1_13, s_1_14, s_1_15, s_1_16, s_1_17, s_1_18, s_1_19, s_1_20, s_1_21, s_1_22, s_1_23, s_1_24, s_1_25, s_1_26, s_1_27, s_1_28, s_1_29, s_1_30, s_1_31, s_1_32;
    wire c_1_1, c_1_2, c_1_3, c_1_4, c_1_5, c_1_6, c_1_7, c_1_8, c_1_9, c_1_10, c_1_11, c_1_12, c_1_13, c_1_14, c_1_15, c_1_16, c_1_17, c_1_18, c_1_19, c_1_20, c_1_21, c_1_22, c_1_23, c_1_24, c_1_25, c_1_26, c_1_27, c_1_28, c_1_29, c_1_30, c_1_31, c_1_32;
    assign w_1_1 = data_operandA[0] & data_operandB[1];
    assign w_1_2 = data_operandA[1] & data_operandB[1];
    assign w_1_3 = data_operandA[2] & data_operandB[1];
    assign w_1_4 = data_operandA[3] & data_operandB[1];
    assign w_1_5 = data_operandA[4] & data_operandB[1];
    assign w_1_6 = data_operandA[5] & data_operandB[1];
    assign w_1_7 = data_operandA[6] & data_operandB[1];
    assign w_1_8 = data_operandA[7] & data_operandB[1];
    assign w_1_9 = data_operandA[8] & data_operandB[1];
    assign w_1_10 = data_operandA[9] & data_operandB[1];
    assign w_1_11 = data_operandA[10] & data_operandB[1];
    assign w_1_12 = data_operandA[11] & data_operandB[1];
    assign w_1_13 = data_operandA[12] & data_operandB[1];
    assign w_1_14 = data_operandA[13] & data_operandB[1];
    assign w_1_15 = data_operandA[14] & data_operandB[1];
    assign w_1_16 = data_operandA[15] & data_operandB[1];
    assign w_1_17 = data_operandA[16] & data_operandB[1];
    assign w_1_18 = data_operandA[17] & data_operandB[1];
    assign w_1_19 = data_operandA[18] & data_operandB[1];
    assign w_1_20 = data_operandA[19] & data_operandB[1];
    assign w_1_21 = data_operandA[20] & data_operandB[1];
    assign w_1_22 = data_operandA[21] & data_operandB[1];
    assign w_1_23 = data_operandA[22] & data_operandB[1];
    assign w_1_24 = data_operandA[23] & data_operandB[1];
    assign w_1_25 = data_operandA[24] & data_operandB[1];
    assign w_1_26 = data_operandA[25] & data_operandB[1];
    assign w_1_27 = data_operandA[26] & data_operandB[1];
    assign w_1_28 = data_operandA[27] & data_operandB[1];
    assign w_1_29 = data_operandA[28] & data_operandB[1];
    assign w_1_30 = data_operandA[29] & data_operandB[1];
    assign w_1_31 = data_operandA[30] & data_operandB[1];
    assign w_1_32 = ~(data_operandA[31] & data_operandB[1]);
    full_adder adder_1_1(.S(s_1_1), .Cout(c_1_1), .A(w_0_1), .B(w_1_1), .Cin(1'b0));
    full_adder adder_1_2(.S(s_1_2), .Cout(c_1_2), .A(w_0_2), .B(w_1_2), .Cin(c_1_1));
    full_adder adder_1_3(.S(s_1_3), .Cout(c_1_3), .A(w_0_3), .B(w_1_3), .Cin(c_1_2));
    full_adder adder_1_4(.S(s_1_4), .Cout(c_1_4), .A(w_0_4), .B(w_1_4), .Cin(c_1_3));
    full_adder adder_1_5(.S(s_1_5), .Cout(c_1_5), .A(w_0_5), .B(w_1_5), .Cin(c_1_4));
    full_adder adder_1_6(.S(s_1_6), .Cout(c_1_6), .A(w_0_6), .B(w_1_6), .Cin(c_1_5));
    full_adder adder_1_7(.S(s_1_7), .Cout(c_1_7), .A(w_0_7), .B(w_1_7), .Cin(c_1_6));
    full_adder adder_1_8(.S(s_1_8), .Cout(c_1_8), .A(w_0_8), .B(w_1_8), .Cin(c_1_7));
    full_adder adder_1_9(.S(s_1_9), .Cout(c_1_9), .A(w_0_9), .B(w_1_9), .Cin(c_1_8));
    full_adder adder_1_10(.S(s_1_10), .Cout(c_1_10), .A(w_0_10), .B(w_1_10), .Cin(c_1_9));
    full_adder adder_1_11(.S(s_1_11), .Cout(c_1_11), .A(w_0_11), .B(w_1_11), .Cin(c_1_10));
    full_adder adder_1_12(.S(s_1_12), .Cout(c_1_12), .A(w_0_12), .B(w_1_12), .Cin(c_1_11));
    full_adder adder_1_13(.S(s_1_13), .Cout(c_1_13), .A(w_0_13), .B(w_1_13), .Cin(c_1_12));
    full_adder adder_1_14(.S(s_1_14), .Cout(c_1_14), .A(w_0_14), .B(w_1_14), .Cin(c_1_13));
    full_adder adder_1_15(.S(s_1_15), .Cout(c_1_15), .A(w_0_15), .B(w_1_15), .Cin(c_1_14));
    full_adder adder_1_16(.S(s_1_16), .Cout(c_1_16), .A(w_0_16), .B(w_1_16), .Cin(c_1_15));
    full_adder adder_1_17(.S(s_1_17), .Cout(c_1_17), .A(w_0_17), .B(w_1_17), .Cin(c_1_16));
    full_adder adder_1_18(.S(s_1_18), .Cout(c_1_18), .A(w_0_18), .B(w_1_18), .Cin(c_1_17));
    full_adder adder_1_19(.S(s_1_19), .Cout(c_1_19), .A(w_0_19), .B(w_1_19), .Cin(c_1_18));
    full_adder adder_1_20(.S(s_1_20), .Cout(c_1_20), .A(w_0_20), .B(w_1_20), .Cin(c_1_19));
    full_adder adder_1_21(.S(s_1_21), .Cout(c_1_21), .A(w_0_21), .B(w_1_21), .Cin(c_1_20));
    full_adder adder_1_22(.S(s_1_22), .Cout(c_1_22), .A(w_0_22), .B(w_1_22), .Cin(c_1_21));
    full_adder adder_1_23(.S(s_1_23), .Cout(c_1_23), .A(w_0_23), .B(w_1_23), .Cin(c_1_22));
    full_adder adder_1_24(.S(s_1_24), .Cout(c_1_24), .A(w_0_24), .B(w_1_24), .Cin(c_1_23));
    full_adder adder_1_25(.S(s_1_25), .Cout(c_1_25), .A(w_0_25), .B(w_1_25), .Cin(c_1_24));
    full_adder adder_1_26(.S(s_1_26), .Cout(c_1_26), .A(w_0_26), .B(w_1_26), .Cin(c_1_25));
    full_adder adder_1_27(.S(s_1_27), .Cout(c_1_27), .A(w_0_27), .B(w_1_27), .Cin(c_1_26));
    full_adder adder_1_28(.S(s_1_28), .Cout(c_1_28), .A(w_0_28), .B(w_1_28), .Cin(c_1_27));
    full_adder adder_1_29(.S(s_1_29), .Cout(c_1_29), .A(w_0_29), .B(w_1_29), .Cin(c_1_28));
    full_adder adder_1_30(.S(s_1_30), .Cout(c_1_30), .A(w_0_30), .B(w_1_30), .Cin(c_1_29));
    full_adder adder_1_31(.S(s_1_31), .Cout(c_1_31), .A(w_0_31), .B(w_1_31), .Cin(c_1_30));
    full_adder adder_1_32(.S(s_1_32), .Cout(c_1_32), .A(1'b1), .B(w_1_32), .Cin(c_1_31));
    assign result[1] = s_1_1;
    wire w_2_2, w_2_3, w_2_4, w_2_5, w_2_6, w_2_7, w_2_8, w_2_9, w_2_10, w_2_11, w_2_12, w_2_13, w_2_14, w_2_15, w_2_16, w_2_17, w_2_18, w_2_19, w_2_20, w_2_21, w_2_22, w_2_23, w_2_24, w_2_25, w_2_26, w_2_27, w_2_28, w_2_29, w_2_30, w_2_31, w_2_32, w_2_33;
    wire s_2_2, s_2_3, s_2_4, s_2_5, s_2_6, s_2_7, s_2_8, s_2_9, s_2_10, s_2_11, s_2_12, s_2_13, s_2_14, s_2_15, s_2_16, s_2_17, s_2_18, s_2_19, s_2_20, s_2_21, s_2_22, s_2_23, s_2_24, s_2_25, s_2_26, s_2_27, s_2_28, s_2_29, s_2_30, s_2_31, s_2_32, s_2_33;
    wire c_2_2, c_2_3, c_2_4, c_2_5, c_2_6, c_2_7, c_2_8, c_2_9, c_2_10, c_2_11, c_2_12, c_2_13, c_2_14, c_2_15, c_2_16, c_2_17, c_2_18, c_2_19, c_2_20, c_2_21, c_2_22, c_2_23, c_2_24, c_2_25, c_2_26, c_2_27, c_2_28, c_2_29, c_2_30, c_2_31, c_2_32, c_2_33;
    assign w_2_2 = data_operandA[0] & data_operandB[2];
    assign w_2_3 = data_operandA[1] & data_operandB[2];
    assign w_2_4 = data_operandA[2] & data_operandB[2];
    assign w_2_5 = data_operandA[3] & data_operandB[2];
    assign w_2_6 = data_operandA[4] & data_operandB[2];
    assign w_2_7 = data_operandA[5] & data_operandB[2];
    assign w_2_8 = data_operandA[6] & data_operandB[2];
    assign w_2_9 = data_operandA[7] & data_operandB[2];
    assign w_2_10 = data_operandA[8] & data_operandB[2];
    assign w_2_11 = data_operandA[9] & data_operandB[2];
    assign w_2_12 = data_operandA[10] & data_operandB[2];
    assign w_2_13 = data_operandA[11] & data_operandB[2];
    assign w_2_14 = data_operandA[12] & data_operandB[2];
    assign w_2_15 = data_operandA[13] & data_operandB[2];
    assign w_2_16 = data_operandA[14] & data_operandB[2];
    assign w_2_17 = data_operandA[15] & data_operandB[2];
    assign w_2_18 = data_operandA[16] & data_operandB[2];
    assign w_2_19 = data_operandA[17] & data_operandB[2];
    assign w_2_20 = data_operandA[18] & data_operandB[2];
    assign w_2_21 = data_operandA[19] & data_operandB[2];
    assign w_2_22 = data_operandA[20] & data_operandB[2];
    assign w_2_23 = data_operandA[21] & data_operandB[2];
    assign w_2_24 = data_operandA[22] & data_operandB[2];
    assign w_2_25 = data_operandA[23] & data_operandB[2];
    assign w_2_26 = data_operandA[24] & data_operandB[2];
    assign w_2_27 = data_operandA[25] & data_operandB[2];
    assign w_2_28 = data_operandA[26] & data_operandB[2];
    assign w_2_29 = data_operandA[27] & data_operandB[2];
    assign w_2_30 = data_operandA[28] & data_operandB[2];
    assign w_2_31 = data_operandA[29] & data_operandB[2];
    assign w_2_32 = data_operandA[30] & data_operandB[2];
    assign w_2_33 = ~(data_operandA[31] & data_operandB[2]);
    full_adder adder_2_2(.S(s_2_2), .Cout(c_2_2), .A(s_1_2), .B(w_2_2), .Cin(1'b0));
    full_adder adder_2_3(.S(s_2_3), .Cout(c_2_3), .A(s_1_3), .B(w_2_3), .Cin(c_2_2));
    full_adder adder_2_4(.S(s_2_4), .Cout(c_2_4), .A(s_1_4), .B(w_2_4), .Cin(c_2_3));
    full_adder adder_2_5(.S(s_2_5), .Cout(c_2_5), .A(s_1_5), .B(w_2_5), .Cin(c_2_4));
    full_adder adder_2_6(.S(s_2_6), .Cout(c_2_6), .A(s_1_6), .B(w_2_6), .Cin(c_2_5));
    full_adder adder_2_7(.S(s_2_7), .Cout(c_2_7), .A(s_1_7), .B(w_2_7), .Cin(c_2_6));
    full_adder adder_2_8(.S(s_2_8), .Cout(c_2_8), .A(s_1_8), .B(w_2_8), .Cin(c_2_7));
    full_adder adder_2_9(.S(s_2_9), .Cout(c_2_9), .A(s_1_9), .B(w_2_9), .Cin(c_2_8));
    full_adder adder_2_10(.S(s_2_10), .Cout(c_2_10), .A(s_1_10), .B(w_2_10), .Cin(c_2_9));
    full_adder adder_2_11(.S(s_2_11), .Cout(c_2_11), .A(s_1_11), .B(w_2_11), .Cin(c_2_10));
    full_adder adder_2_12(.S(s_2_12), .Cout(c_2_12), .A(s_1_12), .B(w_2_12), .Cin(c_2_11));
    full_adder adder_2_13(.S(s_2_13), .Cout(c_2_13), .A(s_1_13), .B(w_2_13), .Cin(c_2_12));
    full_adder adder_2_14(.S(s_2_14), .Cout(c_2_14), .A(s_1_14), .B(w_2_14), .Cin(c_2_13));
    full_adder adder_2_15(.S(s_2_15), .Cout(c_2_15), .A(s_1_15), .B(w_2_15), .Cin(c_2_14));
    full_adder adder_2_16(.S(s_2_16), .Cout(c_2_16), .A(s_1_16), .B(w_2_16), .Cin(c_2_15));
    full_adder adder_2_17(.S(s_2_17), .Cout(c_2_17), .A(s_1_17), .B(w_2_17), .Cin(c_2_16));
    full_adder adder_2_18(.S(s_2_18), .Cout(c_2_18), .A(s_1_18), .B(w_2_18), .Cin(c_2_17));
    full_adder adder_2_19(.S(s_2_19), .Cout(c_2_19), .A(s_1_19), .B(w_2_19), .Cin(c_2_18));
    full_adder adder_2_20(.S(s_2_20), .Cout(c_2_20), .A(s_1_20), .B(w_2_20), .Cin(c_2_19));
    full_adder adder_2_21(.S(s_2_21), .Cout(c_2_21), .A(s_1_21), .B(w_2_21), .Cin(c_2_20));
    full_adder adder_2_22(.S(s_2_22), .Cout(c_2_22), .A(s_1_22), .B(w_2_22), .Cin(c_2_21));
    full_adder adder_2_23(.S(s_2_23), .Cout(c_2_23), .A(s_1_23), .B(w_2_23), .Cin(c_2_22));
    full_adder adder_2_24(.S(s_2_24), .Cout(c_2_24), .A(s_1_24), .B(w_2_24), .Cin(c_2_23));
    full_adder adder_2_25(.S(s_2_25), .Cout(c_2_25), .A(s_1_25), .B(w_2_25), .Cin(c_2_24));
    full_adder adder_2_26(.S(s_2_26), .Cout(c_2_26), .A(s_1_26), .B(w_2_26), .Cin(c_2_25));
    full_adder adder_2_27(.S(s_2_27), .Cout(c_2_27), .A(s_1_27), .B(w_2_27), .Cin(c_2_26));
    full_adder adder_2_28(.S(s_2_28), .Cout(c_2_28), .A(s_1_28), .B(w_2_28), .Cin(c_2_27));
    full_adder adder_2_29(.S(s_2_29), .Cout(c_2_29), .A(s_1_29), .B(w_2_29), .Cin(c_2_28));
    full_adder adder_2_30(.S(s_2_30), .Cout(c_2_30), .A(s_1_30), .B(w_2_30), .Cin(c_2_29));
    full_adder adder_2_31(.S(s_2_31), .Cout(c_2_31), .A(s_1_31), .B(w_2_31), .Cin(c_2_30));
    full_adder adder_2_32(.S(s_2_32), .Cout(c_2_32), .A(s_1_32), .B(w_2_32), .Cin(c_2_31));
    full_adder adder_2_33(.S(s_2_33), .Cout(c_2_33), .A(c_1_32), .B(w_2_33), .Cin(c_2_32));
    assign result[2] = s_2_2;
    wire w_3_3, w_3_4, w_3_5, w_3_6, w_3_7, w_3_8, w_3_9, w_3_10, w_3_11, w_3_12, w_3_13, w_3_14, w_3_15, w_3_16, w_3_17, w_3_18, w_3_19, w_3_20, w_3_21, w_3_22, w_3_23, w_3_24, w_3_25, w_3_26, w_3_27, w_3_28, w_3_29, w_3_30, w_3_31, w_3_32, w_3_33, w_3_34;
    wire s_3_3, s_3_4, s_3_5, s_3_6, s_3_7, s_3_8, s_3_9, s_3_10, s_3_11, s_3_12, s_3_13, s_3_14, s_3_15, s_3_16, s_3_17, s_3_18, s_3_19, s_3_20, s_3_21, s_3_22, s_3_23, s_3_24, s_3_25, s_3_26, s_3_27, s_3_28, s_3_29, s_3_30, s_3_31, s_3_32, s_3_33, s_3_34;
    wire c_3_3, c_3_4, c_3_5, c_3_6, c_3_7, c_3_8, c_3_9, c_3_10, c_3_11, c_3_12, c_3_13, c_3_14, c_3_15, c_3_16, c_3_17, c_3_18, c_3_19, c_3_20, c_3_21, c_3_22, c_3_23, c_3_24, c_3_25, c_3_26, c_3_27, c_3_28, c_3_29, c_3_30, c_3_31, c_3_32, c_3_33, c_3_34;
    assign w_3_3 = data_operandA[0] & data_operandB[3];
    assign w_3_4 = data_operandA[1] & data_operandB[3];
    assign w_3_5 = data_operandA[2] & data_operandB[3];
    assign w_3_6 = data_operandA[3] & data_operandB[3];
    assign w_3_7 = data_operandA[4] & data_operandB[3];
    assign w_3_8 = data_operandA[5] & data_operandB[3];
    assign w_3_9 = data_operandA[6] & data_operandB[3];
    assign w_3_10 = data_operandA[7] & data_operandB[3];
    assign w_3_11 = data_operandA[8] & data_operandB[3];
    assign w_3_12 = data_operandA[9] & data_operandB[3];
    assign w_3_13 = data_operandA[10] & data_operandB[3];
    assign w_3_14 = data_operandA[11] & data_operandB[3];
    assign w_3_15 = data_operandA[12] & data_operandB[3];
    assign w_3_16 = data_operandA[13] & data_operandB[3];
    assign w_3_17 = data_operandA[14] & data_operandB[3];
    assign w_3_18 = data_operandA[15] & data_operandB[3];
    assign w_3_19 = data_operandA[16] & data_operandB[3];
    assign w_3_20 = data_operandA[17] & data_operandB[3];
    assign w_3_21 = data_operandA[18] & data_operandB[3];
    assign w_3_22 = data_operandA[19] & data_operandB[3];
    assign w_3_23 = data_operandA[20] & data_operandB[3];
    assign w_3_24 = data_operandA[21] & data_operandB[3];
    assign w_3_25 = data_operandA[22] & data_operandB[3];
    assign w_3_26 = data_operandA[23] & data_operandB[3];
    assign w_3_27 = data_operandA[24] & data_operandB[3];
    assign w_3_28 = data_operandA[25] & data_operandB[3];
    assign w_3_29 = data_operandA[26] & data_operandB[3];
    assign w_3_30 = data_operandA[27] & data_operandB[3];
    assign w_3_31 = data_operandA[28] & data_operandB[3];
    assign w_3_32 = data_operandA[29] & data_operandB[3];
    assign w_3_33 = data_operandA[30] & data_operandB[3];
    assign w_3_34 = ~(data_operandA[31] & data_operandB[3]);
    full_adder adder_3_3(.S(s_3_3), .Cout(c_3_3), .A(s_2_3), .B(w_3_3), .Cin(1'b0));
    full_adder adder_3_4(.S(s_3_4), .Cout(c_3_4), .A(s_2_4), .B(w_3_4), .Cin(c_3_3));
    full_adder adder_3_5(.S(s_3_5), .Cout(c_3_5), .A(s_2_5), .B(w_3_5), .Cin(c_3_4));
    full_adder adder_3_6(.S(s_3_6), .Cout(c_3_6), .A(s_2_6), .B(w_3_6), .Cin(c_3_5));
    full_adder adder_3_7(.S(s_3_7), .Cout(c_3_7), .A(s_2_7), .B(w_3_7), .Cin(c_3_6));
    full_adder adder_3_8(.S(s_3_8), .Cout(c_3_8), .A(s_2_8), .B(w_3_8), .Cin(c_3_7));
    full_adder adder_3_9(.S(s_3_9), .Cout(c_3_9), .A(s_2_9), .B(w_3_9), .Cin(c_3_8));
    full_adder adder_3_10(.S(s_3_10), .Cout(c_3_10), .A(s_2_10), .B(w_3_10), .Cin(c_3_9));
    full_adder adder_3_11(.S(s_3_11), .Cout(c_3_11), .A(s_2_11), .B(w_3_11), .Cin(c_3_10));
    full_adder adder_3_12(.S(s_3_12), .Cout(c_3_12), .A(s_2_12), .B(w_3_12), .Cin(c_3_11));
    full_adder adder_3_13(.S(s_3_13), .Cout(c_3_13), .A(s_2_13), .B(w_3_13), .Cin(c_3_12));
    full_adder adder_3_14(.S(s_3_14), .Cout(c_3_14), .A(s_2_14), .B(w_3_14), .Cin(c_3_13));
    full_adder adder_3_15(.S(s_3_15), .Cout(c_3_15), .A(s_2_15), .B(w_3_15), .Cin(c_3_14));
    full_adder adder_3_16(.S(s_3_16), .Cout(c_3_16), .A(s_2_16), .B(w_3_16), .Cin(c_3_15));
    full_adder adder_3_17(.S(s_3_17), .Cout(c_3_17), .A(s_2_17), .B(w_3_17), .Cin(c_3_16));
    full_adder adder_3_18(.S(s_3_18), .Cout(c_3_18), .A(s_2_18), .B(w_3_18), .Cin(c_3_17));
    full_adder adder_3_19(.S(s_3_19), .Cout(c_3_19), .A(s_2_19), .B(w_3_19), .Cin(c_3_18));
    full_adder adder_3_20(.S(s_3_20), .Cout(c_3_20), .A(s_2_20), .B(w_3_20), .Cin(c_3_19));
    full_adder adder_3_21(.S(s_3_21), .Cout(c_3_21), .A(s_2_21), .B(w_3_21), .Cin(c_3_20));
    full_adder adder_3_22(.S(s_3_22), .Cout(c_3_22), .A(s_2_22), .B(w_3_22), .Cin(c_3_21));
    full_adder adder_3_23(.S(s_3_23), .Cout(c_3_23), .A(s_2_23), .B(w_3_23), .Cin(c_3_22));
    full_adder adder_3_24(.S(s_3_24), .Cout(c_3_24), .A(s_2_24), .B(w_3_24), .Cin(c_3_23));
    full_adder adder_3_25(.S(s_3_25), .Cout(c_3_25), .A(s_2_25), .B(w_3_25), .Cin(c_3_24));
    full_adder adder_3_26(.S(s_3_26), .Cout(c_3_26), .A(s_2_26), .B(w_3_26), .Cin(c_3_25));
    full_adder adder_3_27(.S(s_3_27), .Cout(c_3_27), .A(s_2_27), .B(w_3_27), .Cin(c_3_26));
    full_adder adder_3_28(.S(s_3_28), .Cout(c_3_28), .A(s_2_28), .B(w_3_28), .Cin(c_3_27));
    full_adder adder_3_29(.S(s_3_29), .Cout(c_3_29), .A(s_2_29), .B(w_3_29), .Cin(c_3_28));
    full_adder adder_3_30(.S(s_3_30), .Cout(c_3_30), .A(s_2_30), .B(w_3_30), .Cin(c_3_29));
    full_adder adder_3_31(.S(s_3_31), .Cout(c_3_31), .A(s_2_31), .B(w_3_31), .Cin(c_3_30));
    full_adder adder_3_32(.S(s_3_32), .Cout(c_3_32), .A(s_2_32), .B(w_3_32), .Cin(c_3_31));
    full_adder adder_3_33(.S(s_3_33), .Cout(c_3_33), .A(s_2_33), .B(w_3_33), .Cin(c_3_32));
    full_adder adder_3_34(.S(s_3_34), .Cout(c_3_34), .A(c_2_33), .B(w_3_34), .Cin(c_3_33));
    assign result[3] = s_3_3;
    wire w_4_4, w_4_5, w_4_6, w_4_7, w_4_8, w_4_9, w_4_10, w_4_11, w_4_12, w_4_13, w_4_14, w_4_15, w_4_16, w_4_17, w_4_18, w_4_19, w_4_20, w_4_21, w_4_22, w_4_23, w_4_24, w_4_25, w_4_26, w_4_27, w_4_28, w_4_29, w_4_30, w_4_31, w_4_32, w_4_33, w_4_34, w_4_35;
    wire s_4_4, s_4_5, s_4_6, s_4_7, s_4_8, s_4_9, s_4_10, s_4_11, s_4_12, s_4_13, s_4_14, s_4_15, s_4_16, s_4_17, s_4_18, s_4_19, s_4_20, s_4_21, s_4_22, s_4_23, s_4_24, s_4_25, s_4_26, s_4_27, s_4_28, s_4_29, s_4_30, s_4_31, s_4_32, s_4_33, s_4_34, s_4_35;
    wire c_4_4, c_4_5, c_4_6, c_4_7, c_4_8, c_4_9, c_4_10, c_4_11, c_4_12, c_4_13, c_4_14, c_4_15, c_4_16, c_4_17, c_4_18, c_4_19, c_4_20, c_4_21, c_4_22, c_4_23, c_4_24, c_4_25, c_4_26, c_4_27, c_4_28, c_4_29, c_4_30, c_4_31, c_4_32, c_4_33, c_4_34, c_4_35;
    assign w_4_4 = data_operandA[0] & data_operandB[4];
    assign w_4_5 = data_operandA[1] & data_operandB[4];
    assign w_4_6 = data_operandA[2] & data_operandB[4];
    assign w_4_7 = data_operandA[3] & data_operandB[4];
    assign w_4_8 = data_operandA[4] & data_operandB[4];
    assign w_4_9 = data_operandA[5] & data_operandB[4];
    assign w_4_10 = data_operandA[6] & data_operandB[4];
    assign w_4_11 = data_operandA[7] & data_operandB[4];
    assign w_4_12 = data_operandA[8] & data_operandB[4];
    assign w_4_13 = data_operandA[9] & data_operandB[4];
    assign w_4_14 = data_operandA[10] & data_operandB[4];
    assign w_4_15 = data_operandA[11] & data_operandB[4];
    assign w_4_16 = data_operandA[12] & data_operandB[4];
    assign w_4_17 = data_operandA[13] & data_operandB[4];
    assign w_4_18 = data_operandA[14] & data_operandB[4];
    assign w_4_19 = data_operandA[15] & data_operandB[4];
    assign w_4_20 = data_operandA[16] & data_operandB[4];
    assign w_4_21 = data_operandA[17] & data_operandB[4];
    assign w_4_22 = data_operandA[18] & data_operandB[4];
    assign w_4_23 = data_operandA[19] & data_operandB[4];
    assign w_4_24 = data_operandA[20] & data_operandB[4];
    assign w_4_25 = data_operandA[21] & data_operandB[4];
    assign w_4_26 = data_operandA[22] & data_operandB[4];
    assign w_4_27 = data_operandA[23] & data_operandB[4];
    assign w_4_28 = data_operandA[24] & data_operandB[4];
    assign w_4_29 = data_operandA[25] & data_operandB[4];
    assign w_4_30 = data_operandA[26] & data_operandB[4];
    assign w_4_31 = data_operandA[27] & data_operandB[4];
    assign w_4_32 = data_operandA[28] & data_operandB[4];
    assign w_4_33 = data_operandA[29] & data_operandB[4];
    assign w_4_34 = data_operandA[30] & data_operandB[4];
    assign w_4_35 = ~(data_operandA[31] & data_operandB[4]);
    full_adder adder_4_4(.S(s_4_4), .Cout(c_4_4), .A(s_3_4), .B(w_4_4), .Cin(1'b0));
    full_adder adder_4_5(.S(s_4_5), .Cout(c_4_5), .A(s_3_5), .B(w_4_5), .Cin(c_4_4));
    full_adder adder_4_6(.S(s_4_6), .Cout(c_4_6), .A(s_3_6), .B(w_4_6), .Cin(c_4_5));
    full_adder adder_4_7(.S(s_4_7), .Cout(c_4_7), .A(s_3_7), .B(w_4_7), .Cin(c_4_6));
    full_adder adder_4_8(.S(s_4_8), .Cout(c_4_8), .A(s_3_8), .B(w_4_8), .Cin(c_4_7));
    full_adder adder_4_9(.S(s_4_9), .Cout(c_4_9), .A(s_3_9), .B(w_4_9), .Cin(c_4_8));
    full_adder adder_4_10(.S(s_4_10), .Cout(c_4_10), .A(s_3_10), .B(w_4_10), .Cin(c_4_9));
    full_adder adder_4_11(.S(s_4_11), .Cout(c_4_11), .A(s_3_11), .B(w_4_11), .Cin(c_4_10));
    full_adder adder_4_12(.S(s_4_12), .Cout(c_4_12), .A(s_3_12), .B(w_4_12), .Cin(c_4_11));
    full_adder adder_4_13(.S(s_4_13), .Cout(c_4_13), .A(s_3_13), .B(w_4_13), .Cin(c_4_12));
    full_adder adder_4_14(.S(s_4_14), .Cout(c_4_14), .A(s_3_14), .B(w_4_14), .Cin(c_4_13));
    full_adder adder_4_15(.S(s_4_15), .Cout(c_4_15), .A(s_3_15), .B(w_4_15), .Cin(c_4_14));
    full_adder adder_4_16(.S(s_4_16), .Cout(c_4_16), .A(s_3_16), .B(w_4_16), .Cin(c_4_15));
    full_adder adder_4_17(.S(s_4_17), .Cout(c_4_17), .A(s_3_17), .B(w_4_17), .Cin(c_4_16));
    full_adder adder_4_18(.S(s_4_18), .Cout(c_4_18), .A(s_3_18), .B(w_4_18), .Cin(c_4_17));
    full_adder adder_4_19(.S(s_4_19), .Cout(c_4_19), .A(s_3_19), .B(w_4_19), .Cin(c_4_18));
    full_adder adder_4_20(.S(s_4_20), .Cout(c_4_20), .A(s_3_20), .B(w_4_20), .Cin(c_4_19));
    full_adder adder_4_21(.S(s_4_21), .Cout(c_4_21), .A(s_3_21), .B(w_4_21), .Cin(c_4_20));
    full_adder adder_4_22(.S(s_4_22), .Cout(c_4_22), .A(s_3_22), .B(w_4_22), .Cin(c_4_21));
    full_adder adder_4_23(.S(s_4_23), .Cout(c_4_23), .A(s_3_23), .B(w_4_23), .Cin(c_4_22));
    full_adder adder_4_24(.S(s_4_24), .Cout(c_4_24), .A(s_3_24), .B(w_4_24), .Cin(c_4_23));
    full_adder adder_4_25(.S(s_4_25), .Cout(c_4_25), .A(s_3_25), .B(w_4_25), .Cin(c_4_24));
    full_adder adder_4_26(.S(s_4_26), .Cout(c_4_26), .A(s_3_26), .B(w_4_26), .Cin(c_4_25));
    full_adder adder_4_27(.S(s_4_27), .Cout(c_4_27), .A(s_3_27), .B(w_4_27), .Cin(c_4_26));
    full_adder adder_4_28(.S(s_4_28), .Cout(c_4_28), .A(s_3_28), .B(w_4_28), .Cin(c_4_27));
    full_adder adder_4_29(.S(s_4_29), .Cout(c_4_29), .A(s_3_29), .B(w_4_29), .Cin(c_4_28));
    full_adder adder_4_30(.S(s_4_30), .Cout(c_4_30), .A(s_3_30), .B(w_4_30), .Cin(c_4_29));
    full_adder adder_4_31(.S(s_4_31), .Cout(c_4_31), .A(s_3_31), .B(w_4_31), .Cin(c_4_30));
    full_adder adder_4_32(.S(s_4_32), .Cout(c_4_32), .A(s_3_32), .B(w_4_32), .Cin(c_4_31));
    full_adder adder_4_33(.S(s_4_33), .Cout(c_4_33), .A(s_3_33), .B(w_4_33), .Cin(c_4_32));
    full_adder adder_4_34(.S(s_4_34), .Cout(c_4_34), .A(s_3_34), .B(w_4_34), .Cin(c_4_33));
    full_adder adder_4_35(.S(s_4_35), .Cout(c_4_35), .A(c_3_34), .B(w_4_35), .Cin(c_4_34));
    assign result[4] = s_4_4;
    wire w_5_5, w_5_6, w_5_7, w_5_8, w_5_9, w_5_10, w_5_11, w_5_12, w_5_13, w_5_14, w_5_15, w_5_16, w_5_17, w_5_18, w_5_19, w_5_20, w_5_21, w_5_22, w_5_23, w_5_24, w_5_25, w_5_26, w_5_27, w_5_28, w_5_29, w_5_30, w_5_31, w_5_32, w_5_33, w_5_34, w_5_35, w_5_36;
    wire s_5_5, s_5_6, s_5_7, s_5_8, s_5_9, s_5_10, s_5_11, s_5_12, s_5_13, s_5_14, s_5_15, s_5_16, s_5_17, s_5_18, s_5_19, s_5_20, s_5_21, s_5_22, s_5_23, s_5_24, s_5_25, s_5_26, s_5_27, s_5_28, s_5_29, s_5_30, s_5_31, s_5_32, s_5_33, s_5_34, s_5_35, s_5_36;
    wire c_5_5, c_5_6, c_5_7, c_5_8, c_5_9, c_5_10, c_5_11, c_5_12, c_5_13, c_5_14, c_5_15, c_5_16, c_5_17, c_5_18, c_5_19, c_5_20, c_5_21, c_5_22, c_5_23, c_5_24, c_5_25, c_5_26, c_5_27, c_5_28, c_5_29, c_5_30, c_5_31, c_5_32, c_5_33, c_5_34, c_5_35, c_5_36;
    assign w_5_5 = data_operandA[0] & data_operandB[5];
    assign w_5_6 = data_operandA[1] & data_operandB[5];
    assign w_5_7 = data_operandA[2] & data_operandB[5];
    assign w_5_8 = data_operandA[3] & data_operandB[5];
    assign w_5_9 = data_operandA[4] & data_operandB[5];
    assign w_5_10 = data_operandA[5] & data_operandB[5];
    assign w_5_11 = data_operandA[6] & data_operandB[5];
    assign w_5_12 = data_operandA[7] & data_operandB[5];
    assign w_5_13 = data_operandA[8] & data_operandB[5];
    assign w_5_14 = data_operandA[9] & data_operandB[5];
    assign w_5_15 = data_operandA[10] & data_operandB[5];
    assign w_5_16 = data_operandA[11] & data_operandB[5];
    assign w_5_17 = data_operandA[12] & data_operandB[5];
    assign w_5_18 = data_operandA[13] & data_operandB[5];
    assign w_5_19 = data_operandA[14] & data_operandB[5];
    assign w_5_20 = data_operandA[15] & data_operandB[5];
    assign w_5_21 = data_operandA[16] & data_operandB[5];
    assign w_5_22 = data_operandA[17] & data_operandB[5];
    assign w_5_23 = data_operandA[18] & data_operandB[5];
    assign w_5_24 = data_operandA[19] & data_operandB[5];
    assign w_5_25 = data_operandA[20] & data_operandB[5];
    assign w_5_26 = data_operandA[21] & data_operandB[5];
    assign w_5_27 = data_operandA[22] & data_operandB[5];
    assign w_5_28 = data_operandA[23] & data_operandB[5];
    assign w_5_29 = data_operandA[24] & data_operandB[5];
    assign w_5_30 = data_operandA[25] & data_operandB[5];
    assign w_5_31 = data_operandA[26] & data_operandB[5];
    assign w_5_32 = data_operandA[27] & data_operandB[5];
    assign w_5_33 = data_operandA[28] & data_operandB[5];
    assign w_5_34 = data_operandA[29] & data_operandB[5];
    assign w_5_35 = data_operandA[30] & data_operandB[5];
    assign w_5_36 = ~(data_operandA[31] & data_operandB[5]);
    full_adder adder_5_5(.S(s_5_5), .Cout(c_5_5), .A(s_4_5), .B(w_5_5), .Cin(1'b0));
    full_adder adder_5_6(.S(s_5_6), .Cout(c_5_6), .A(s_4_6), .B(w_5_6), .Cin(c_5_5));
    full_adder adder_5_7(.S(s_5_7), .Cout(c_5_7), .A(s_4_7), .B(w_5_7), .Cin(c_5_6));
    full_adder adder_5_8(.S(s_5_8), .Cout(c_5_8), .A(s_4_8), .B(w_5_8), .Cin(c_5_7));
    full_adder adder_5_9(.S(s_5_9), .Cout(c_5_9), .A(s_4_9), .B(w_5_9), .Cin(c_5_8));
    full_adder adder_5_10(.S(s_5_10), .Cout(c_5_10), .A(s_4_10), .B(w_5_10), .Cin(c_5_9));
    full_adder adder_5_11(.S(s_5_11), .Cout(c_5_11), .A(s_4_11), .B(w_5_11), .Cin(c_5_10));
    full_adder adder_5_12(.S(s_5_12), .Cout(c_5_12), .A(s_4_12), .B(w_5_12), .Cin(c_5_11));
    full_adder adder_5_13(.S(s_5_13), .Cout(c_5_13), .A(s_4_13), .B(w_5_13), .Cin(c_5_12));
    full_adder adder_5_14(.S(s_5_14), .Cout(c_5_14), .A(s_4_14), .B(w_5_14), .Cin(c_5_13));
    full_adder adder_5_15(.S(s_5_15), .Cout(c_5_15), .A(s_4_15), .B(w_5_15), .Cin(c_5_14));
    full_adder adder_5_16(.S(s_5_16), .Cout(c_5_16), .A(s_4_16), .B(w_5_16), .Cin(c_5_15));
    full_adder adder_5_17(.S(s_5_17), .Cout(c_5_17), .A(s_4_17), .B(w_5_17), .Cin(c_5_16));
    full_adder adder_5_18(.S(s_5_18), .Cout(c_5_18), .A(s_4_18), .B(w_5_18), .Cin(c_5_17));
    full_adder adder_5_19(.S(s_5_19), .Cout(c_5_19), .A(s_4_19), .B(w_5_19), .Cin(c_5_18));
    full_adder adder_5_20(.S(s_5_20), .Cout(c_5_20), .A(s_4_20), .B(w_5_20), .Cin(c_5_19));
    full_adder adder_5_21(.S(s_5_21), .Cout(c_5_21), .A(s_4_21), .B(w_5_21), .Cin(c_5_20));
    full_adder adder_5_22(.S(s_5_22), .Cout(c_5_22), .A(s_4_22), .B(w_5_22), .Cin(c_5_21));
    full_adder adder_5_23(.S(s_5_23), .Cout(c_5_23), .A(s_4_23), .B(w_5_23), .Cin(c_5_22));
    full_adder adder_5_24(.S(s_5_24), .Cout(c_5_24), .A(s_4_24), .B(w_5_24), .Cin(c_5_23));
    full_adder adder_5_25(.S(s_5_25), .Cout(c_5_25), .A(s_4_25), .B(w_5_25), .Cin(c_5_24));
    full_adder adder_5_26(.S(s_5_26), .Cout(c_5_26), .A(s_4_26), .B(w_5_26), .Cin(c_5_25));
    full_adder adder_5_27(.S(s_5_27), .Cout(c_5_27), .A(s_4_27), .B(w_5_27), .Cin(c_5_26));
    full_adder adder_5_28(.S(s_5_28), .Cout(c_5_28), .A(s_4_28), .B(w_5_28), .Cin(c_5_27));
    full_adder adder_5_29(.S(s_5_29), .Cout(c_5_29), .A(s_4_29), .B(w_5_29), .Cin(c_5_28));
    full_adder adder_5_30(.S(s_5_30), .Cout(c_5_30), .A(s_4_30), .B(w_5_30), .Cin(c_5_29));
    full_adder adder_5_31(.S(s_5_31), .Cout(c_5_31), .A(s_4_31), .B(w_5_31), .Cin(c_5_30));
    full_adder adder_5_32(.S(s_5_32), .Cout(c_5_32), .A(s_4_32), .B(w_5_32), .Cin(c_5_31));
    full_adder adder_5_33(.S(s_5_33), .Cout(c_5_33), .A(s_4_33), .B(w_5_33), .Cin(c_5_32));
    full_adder adder_5_34(.S(s_5_34), .Cout(c_5_34), .A(s_4_34), .B(w_5_34), .Cin(c_5_33));
    full_adder adder_5_35(.S(s_5_35), .Cout(c_5_35), .A(s_4_35), .B(w_5_35), .Cin(c_5_34));
    full_adder adder_5_36(.S(s_5_36), .Cout(c_5_36), .A(c_4_35), .B(w_5_36), .Cin(c_5_35));
    assign result[5] = s_5_5;
    wire w_6_6, w_6_7, w_6_8, w_6_9, w_6_10, w_6_11, w_6_12, w_6_13, w_6_14, w_6_15, w_6_16, w_6_17, w_6_18, w_6_19, w_6_20, w_6_21, w_6_22, w_6_23, w_6_24, w_6_25, w_6_26, w_6_27, w_6_28, w_6_29, w_6_30, w_6_31, w_6_32, w_6_33, w_6_34, w_6_35, w_6_36, w_6_37;
    wire s_6_6, s_6_7, s_6_8, s_6_9, s_6_10, s_6_11, s_6_12, s_6_13, s_6_14, s_6_15, s_6_16, s_6_17, s_6_18, s_6_19, s_6_20, s_6_21, s_6_22, s_6_23, s_6_24, s_6_25, s_6_26, s_6_27, s_6_28, s_6_29, s_6_30, s_6_31, s_6_32, s_6_33, s_6_34, s_6_35, s_6_36, s_6_37;
    wire c_6_6, c_6_7, c_6_8, c_6_9, c_6_10, c_6_11, c_6_12, c_6_13, c_6_14, c_6_15, c_6_16, c_6_17, c_6_18, c_6_19, c_6_20, c_6_21, c_6_22, c_6_23, c_6_24, c_6_25, c_6_26, c_6_27, c_6_28, c_6_29, c_6_30, c_6_31, c_6_32, c_6_33, c_6_34, c_6_35, c_6_36, c_6_37;
    assign w_6_6 = data_operandA[0] & data_operandB[6];
    assign w_6_7 = data_operandA[1] & data_operandB[6];
    assign w_6_8 = data_operandA[2] & data_operandB[6];
    assign w_6_9 = data_operandA[3] & data_operandB[6];
    assign w_6_10 = data_operandA[4] & data_operandB[6];
    assign w_6_11 = data_operandA[5] & data_operandB[6];
    assign w_6_12 = data_operandA[6] & data_operandB[6];
    assign w_6_13 = data_operandA[7] & data_operandB[6];
    assign w_6_14 = data_operandA[8] & data_operandB[6];
    assign w_6_15 = data_operandA[9] & data_operandB[6];
    assign w_6_16 = data_operandA[10] & data_operandB[6];
    assign w_6_17 = data_operandA[11] & data_operandB[6];
    assign w_6_18 = data_operandA[12] & data_operandB[6];
    assign w_6_19 = data_operandA[13] & data_operandB[6];
    assign w_6_20 = data_operandA[14] & data_operandB[6];
    assign w_6_21 = data_operandA[15] & data_operandB[6];
    assign w_6_22 = data_operandA[16] & data_operandB[6];
    assign w_6_23 = data_operandA[17] & data_operandB[6];
    assign w_6_24 = data_operandA[18] & data_operandB[6];
    assign w_6_25 = data_operandA[19] & data_operandB[6];
    assign w_6_26 = data_operandA[20] & data_operandB[6];
    assign w_6_27 = data_operandA[21] & data_operandB[6];
    assign w_6_28 = data_operandA[22] & data_operandB[6];
    assign w_6_29 = data_operandA[23] & data_operandB[6];
    assign w_6_30 = data_operandA[24] & data_operandB[6];
    assign w_6_31 = data_operandA[25] & data_operandB[6];
    assign w_6_32 = data_operandA[26] & data_operandB[6];
    assign w_6_33 = data_operandA[27] & data_operandB[6];
    assign w_6_34 = data_operandA[28] & data_operandB[6];
    assign w_6_35 = data_operandA[29] & data_operandB[6];
    assign w_6_36 = data_operandA[30] & data_operandB[6];
    assign w_6_37 = ~(data_operandA[31] & data_operandB[6]);
    full_adder adder_6_6(.S(s_6_6), .Cout(c_6_6), .A(s_5_6), .B(w_6_6), .Cin(1'b0));
    full_adder adder_6_7(.S(s_6_7), .Cout(c_6_7), .A(s_5_7), .B(w_6_7), .Cin(c_6_6));
    full_adder adder_6_8(.S(s_6_8), .Cout(c_6_8), .A(s_5_8), .B(w_6_8), .Cin(c_6_7));
    full_adder adder_6_9(.S(s_6_9), .Cout(c_6_9), .A(s_5_9), .B(w_6_9), .Cin(c_6_8));
    full_adder adder_6_10(.S(s_6_10), .Cout(c_6_10), .A(s_5_10), .B(w_6_10), .Cin(c_6_9));
    full_adder adder_6_11(.S(s_6_11), .Cout(c_6_11), .A(s_5_11), .B(w_6_11), .Cin(c_6_10));
    full_adder adder_6_12(.S(s_6_12), .Cout(c_6_12), .A(s_5_12), .B(w_6_12), .Cin(c_6_11));
    full_adder adder_6_13(.S(s_6_13), .Cout(c_6_13), .A(s_5_13), .B(w_6_13), .Cin(c_6_12));
    full_adder adder_6_14(.S(s_6_14), .Cout(c_6_14), .A(s_5_14), .B(w_6_14), .Cin(c_6_13));
    full_adder adder_6_15(.S(s_6_15), .Cout(c_6_15), .A(s_5_15), .B(w_6_15), .Cin(c_6_14));
    full_adder adder_6_16(.S(s_6_16), .Cout(c_6_16), .A(s_5_16), .B(w_6_16), .Cin(c_6_15));
    full_adder adder_6_17(.S(s_6_17), .Cout(c_6_17), .A(s_5_17), .B(w_6_17), .Cin(c_6_16));
    full_adder adder_6_18(.S(s_6_18), .Cout(c_6_18), .A(s_5_18), .B(w_6_18), .Cin(c_6_17));
    full_adder adder_6_19(.S(s_6_19), .Cout(c_6_19), .A(s_5_19), .B(w_6_19), .Cin(c_6_18));
    full_adder adder_6_20(.S(s_6_20), .Cout(c_6_20), .A(s_5_20), .B(w_6_20), .Cin(c_6_19));
    full_adder adder_6_21(.S(s_6_21), .Cout(c_6_21), .A(s_5_21), .B(w_6_21), .Cin(c_6_20));
    full_adder adder_6_22(.S(s_6_22), .Cout(c_6_22), .A(s_5_22), .B(w_6_22), .Cin(c_6_21));
    full_adder adder_6_23(.S(s_6_23), .Cout(c_6_23), .A(s_5_23), .B(w_6_23), .Cin(c_6_22));
    full_adder adder_6_24(.S(s_6_24), .Cout(c_6_24), .A(s_5_24), .B(w_6_24), .Cin(c_6_23));
    full_adder adder_6_25(.S(s_6_25), .Cout(c_6_25), .A(s_5_25), .B(w_6_25), .Cin(c_6_24));
    full_adder adder_6_26(.S(s_6_26), .Cout(c_6_26), .A(s_5_26), .B(w_6_26), .Cin(c_6_25));
    full_adder adder_6_27(.S(s_6_27), .Cout(c_6_27), .A(s_5_27), .B(w_6_27), .Cin(c_6_26));
    full_adder adder_6_28(.S(s_6_28), .Cout(c_6_28), .A(s_5_28), .B(w_6_28), .Cin(c_6_27));
    full_adder adder_6_29(.S(s_6_29), .Cout(c_6_29), .A(s_5_29), .B(w_6_29), .Cin(c_6_28));
    full_adder adder_6_30(.S(s_6_30), .Cout(c_6_30), .A(s_5_30), .B(w_6_30), .Cin(c_6_29));
    full_adder adder_6_31(.S(s_6_31), .Cout(c_6_31), .A(s_5_31), .B(w_6_31), .Cin(c_6_30));
    full_adder adder_6_32(.S(s_6_32), .Cout(c_6_32), .A(s_5_32), .B(w_6_32), .Cin(c_6_31));
    full_adder adder_6_33(.S(s_6_33), .Cout(c_6_33), .A(s_5_33), .B(w_6_33), .Cin(c_6_32));
    full_adder adder_6_34(.S(s_6_34), .Cout(c_6_34), .A(s_5_34), .B(w_6_34), .Cin(c_6_33));
    full_adder adder_6_35(.S(s_6_35), .Cout(c_6_35), .A(s_5_35), .B(w_6_35), .Cin(c_6_34));
    full_adder adder_6_36(.S(s_6_36), .Cout(c_6_36), .A(s_5_36), .B(w_6_36), .Cin(c_6_35));
    full_adder adder_6_37(.S(s_6_37), .Cout(c_6_37), .A(c_5_36), .B(w_6_37), .Cin(c_6_36));
    assign result[6] = s_6_6;
    wire w_7_7, w_7_8, w_7_9, w_7_10, w_7_11, w_7_12, w_7_13, w_7_14, w_7_15, w_7_16, w_7_17, w_7_18, w_7_19, w_7_20, w_7_21, w_7_22, w_7_23, w_7_24, w_7_25, w_7_26, w_7_27, w_7_28, w_7_29, w_7_30, w_7_31, w_7_32, w_7_33, w_7_34, w_7_35, w_7_36, w_7_37, w_7_38;
    wire s_7_7, s_7_8, s_7_9, s_7_10, s_7_11, s_7_12, s_7_13, s_7_14, s_7_15, s_7_16, s_7_17, s_7_18, s_7_19, s_7_20, s_7_21, s_7_22, s_7_23, s_7_24, s_7_25, s_7_26, s_7_27, s_7_28, s_7_29, s_7_30, s_7_31, s_7_32, s_7_33, s_7_34, s_7_35, s_7_36, s_7_37, s_7_38;
    wire c_7_7, c_7_8, c_7_9, c_7_10, c_7_11, c_7_12, c_7_13, c_7_14, c_7_15, c_7_16, c_7_17, c_7_18, c_7_19, c_7_20, c_7_21, c_7_22, c_7_23, c_7_24, c_7_25, c_7_26, c_7_27, c_7_28, c_7_29, c_7_30, c_7_31, c_7_32, c_7_33, c_7_34, c_7_35, c_7_36, c_7_37, c_7_38;
    assign w_7_7 = data_operandA[0] & data_operandB[7];
    assign w_7_8 = data_operandA[1] & data_operandB[7];
    assign w_7_9 = data_operandA[2] & data_operandB[7];
    assign w_7_10 = data_operandA[3] & data_operandB[7];
    assign w_7_11 = data_operandA[4] & data_operandB[7];
    assign w_7_12 = data_operandA[5] & data_operandB[7];
    assign w_7_13 = data_operandA[6] & data_operandB[7];
    assign w_7_14 = data_operandA[7] & data_operandB[7];
    assign w_7_15 = data_operandA[8] & data_operandB[7];
    assign w_7_16 = data_operandA[9] & data_operandB[7];
    assign w_7_17 = data_operandA[10] & data_operandB[7];
    assign w_7_18 = data_operandA[11] & data_operandB[7];
    assign w_7_19 = data_operandA[12] & data_operandB[7];
    assign w_7_20 = data_operandA[13] & data_operandB[7];
    assign w_7_21 = data_operandA[14] & data_operandB[7];
    assign w_7_22 = data_operandA[15] & data_operandB[7];
    assign w_7_23 = data_operandA[16] & data_operandB[7];
    assign w_7_24 = data_operandA[17] & data_operandB[7];
    assign w_7_25 = data_operandA[18] & data_operandB[7];
    assign w_7_26 = data_operandA[19] & data_operandB[7];
    assign w_7_27 = data_operandA[20] & data_operandB[7];
    assign w_7_28 = data_operandA[21] & data_operandB[7];
    assign w_7_29 = data_operandA[22] & data_operandB[7];
    assign w_7_30 = data_operandA[23] & data_operandB[7];
    assign w_7_31 = data_operandA[24] & data_operandB[7];
    assign w_7_32 = data_operandA[25] & data_operandB[7];
    assign w_7_33 = data_operandA[26] & data_operandB[7];
    assign w_7_34 = data_operandA[27] & data_operandB[7];
    assign w_7_35 = data_operandA[28] & data_operandB[7];
    assign w_7_36 = data_operandA[29] & data_operandB[7];
    assign w_7_37 = data_operandA[30] & data_operandB[7];
    assign w_7_38 = ~(data_operandA[31] & data_operandB[7]);
    full_adder adder_7_7(.S(s_7_7), .Cout(c_7_7), .A(s_6_7), .B(w_7_7), .Cin(1'b0));
    full_adder adder_7_8(.S(s_7_8), .Cout(c_7_8), .A(s_6_8), .B(w_7_8), .Cin(c_7_7));
    full_adder adder_7_9(.S(s_7_9), .Cout(c_7_9), .A(s_6_9), .B(w_7_9), .Cin(c_7_8));
    full_adder adder_7_10(.S(s_7_10), .Cout(c_7_10), .A(s_6_10), .B(w_7_10), .Cin(c_7_9));
    full_adder adder_7_11(.S(s_7_11), .Cout(c_7_11), .A(s_6_11), .B(w_7_11), .Cin(c_7_10));
    full_adder adder_7_12(.S(s_7_12), .Cout(c_7_12), .A(s_6_12), .B(w_7_12), .Cin(c_7_11));
    full_adder adder_7_13(.S(s_7_13), .Cout(c_7_13), .A(s_6_13), .B(w_7_13), .Cin(c_7_12));
    full_adder adder_7_14(.S(s_7_14), .Cout(c_7_14), .A(s_6_14), .B(w_7_14), .Cin(c_7_13));
    full_adder adder_7_15(.S(s_7_15), .Cout(c_7_15), .A(s_6_15), .B(w_7_15), .Cin(c_7_14));
    full_adder adder_7_16(.S(s_7_16), .Cout(c_7_16), .A(s_6_16), .B(w_7_16), .Cin(c_7_15));
    full_adder adder_7_17(.S(s_7_17), .Cout(c_7_17), .A(s_6_17), .B(w_7_17), .Cin(c_7_16));
    full_adder adder_7_18(.S(s_7_18), .Cout(c_7_18), .A(s_6_18), .B(w_7_18), .Cin(c_7_17));
    full_adder adder_7_19(.S(s_7_19), .Cout(c_7_19), .A(s_6_19), .B(w_7_19), .Cin(c_7_18));
    full_adder adder_7_20(.S(s_7_20), .Cout(c_7_20), .A(s_6_20), .B(w_7_20), .Cin(c_7_19));
    full_adder adder_7_21(.S(s_7_21), .Cout(c_7_21), .A(s_6_21), .B(w_7_21), .Cin(c_7_20));
    full_adder adder_7_22(.S(s_7_22), .Cout(c_7_22), .A(s_6_22), .B(w_7_22), .Cin(c_7_21));
    full_adder adder_7_23(.S(s_7_23), .Cout(c_7_23), .A(s_6_23), .B(w_7_23), .Cin(c_7_22));
    full_adder adder_7_24(.S(s_7_24), .Cout(c_7_24), .A(s_6_24), .B(w_7_24), .Cin(c_7_23));
    full_adder adder_7_25(.S(s_7_25), .Cout(c_7_25), .A(s_6_25), .B(w_7_25), .Cin(c_7_24));
    full_adder adder_7_26(.S(s_7_26), .Cout(c_7_26), .A(s_6_26), .B(w_7_26), .Cin(c_7_25));
    full_adder adder_7_27(.S(s_7_27), .Cout(c_7_27), .A(s_6_27), .B(w_7_27), .Cin(c_7_26));
    full_adder adder_7_28(.S(s_7_28), .Cout(c_7_28), .A(s_6_28), .B(w_7_28), .Cin(c_7_27));
    full_adder adder_7_29(.S(s_7_29), .Cout(c_7_29), .A(s_6_29), .B(w_7_29), .Cin(c_7_28));
    full_adder adder_7_30(.S(s_7_30), .Cout(c_7_30), .A(s_6_30), .B(w_7_30), .Cin(c_7_29));
    full_adder adder_7_31(.S(s_7_31), .Cout(c_7_31), .A(s_6_31), .B(w_7_31), .Cin(c_7_30));
    full_adder adder_7_32(.S(s_7_32), .Cout(c_7_32), .A(s_6_32), .B(w_7_32), .Cin(c_7_31));
    full_adder adder_7_33(.S(s_7_33), .Cout(c_7_33), .A(s_6_33), .B(w_7_33), .Cin(c_7_32));
    full_adder adder_7_34(.S(s_7_34), .Cout(c_7_34), .A(s_6_34), .B(w_7_34), .Cin(c_7_33));
    full_adder adder_7_35(.S(s_7_35), .Cout(c_7_35), .A(s_6_35), .B(w_7_35), .Cin(c_7_34));
    full_adder adder_7_36(.S(s_7_36), .Cout(c_7_36), .A(s_6_36), .B(w_7_36), .Cin(c_7_35));
    full_adder adder_7_37(.S(s_7_37), .Cout(c_7_37), .A(s_6_37), .B(w_7_37), .Cin(c_7_36));
    full_adder adder_7_38(.S(s_7_38), .Cout(c_7_38), .A(c_6_37), .B(w_7_38), .Cin(c_7_37));
    assign result[7] = s_7_7;
    wire w_8_8, w_8_9, w_8_10, w_8_11, w_8_12, w_8_13, w_8_14, w_8_15, w_8_16, w_8_17, w_8_18, w_8_19, w_8_20, w_8_21, w_8_22, w_8_23, w_8_24, w_8_25, w_8_26, w_8_27, w_8_28, w_8_29, w_8_30, w_8_31, w_8_32, w_8_33, w_8_34, w_8_35, w_8_36, w_8_37, w_8_38, w_8_39;
    wire s_8_8, s_8_9, s_8_10, s_8_11, s_8_12, s_8_13, s_8_14, s_8_15, s_8_16, s_8_17, s_8_18, s_8_19, s_8_20, s_8_21, s_8_22, s_8_23, s_8_24, s_8_25, s_8_26, s_8_27, s_8_28, s_8_29, s_8_30, s_8_31, s_8_32, s_8_33, s_8_34, s_8_35, s_8_36, s_8_37, s_8_38, s_8_39;
    wire c_8_8, c_8_9, c_8_10, c_8_11, c_8_12, c_8_13, c_8_14, c_8_15, c_8_16, c_8_17, c_8_18, c_8_19, c_8_20, c_8_21, c_8_22, c_8_23, c_8_24, c_8_25, c_8_26, c_8_27, c_8_28, c_8_29, c_8_30, c_8_31, c_8_32, c_8_33, c_8_34, c_8_35, c_8_36, c_8_37, c_8_38, c_8_39;
    assign w_8_8 = data_operandA[0] & data_operandB[8];
    assign w_8_9 = data_operandA[1] & data_operandB[8];
    assign w_8_10 = data_operandA[2] & data_operandB[8];
    assign w_8_11 = data_operandA[3] & data_operandB[8];
    assign w_8_12 = data_operandA[4] & data_operandB[8];
    assign w_8_13 = data_operandA[5] & data_operandB[8];
    assign w_8_14 = data_operandA[6] & data_operandB[8];
    assign w_8_15 = data_operandA[7] & data_operandB[8];
    assign w_8_16 = data_operandA[8] & data_operandB[8];
    assign w_8_17 = data_operandA[9] & data_operandB[8];
    assign w_8_18 = data_operandA[10] & data_operandB[8];
    assign w_8_19 = data_operandA[11] & data_operandB[8];
    assign w_8_20 = data_operandA[12] & data_operandB[8];
    assign w_8_21 = data_operandA[13] & data_operandB[8];
    assign w_8_22 = data_operandA[14] & data_operandB[8];
    assign w_8_23 = data_operandA[15] & data_operandB[8];
    assign w_8_24 = data_operandA[16] & data_operandB[8];
    assign w_8_25 = data_operandA[17] & data_operandB[8];
    assign w_8_26 = data_operandA[18] & data_operandB[8];
    assign w_8_27 = data_operandA[19] & data_operandB[8];
    assign w_8_28 = data_operandA[20] & data_operandB[8];
    assign w_8_29 = data_operandA[21] & data_operandB[8];
    assign w_8_30 = data_operandA[22] & data_operandB[8];
    assign w_8_31 = data_operandA[23] & data_operandB[8];
    assign w_8_32 = data_operandA[24] & data_operandB[8];
    assign w_8_33 = data_operandA[25] & data_operandB[8];
    assign w_8_34 = data_operandA[26] & data_operandB[8];
    assign w_8_35 = data_operandA[27] & data_operandB[8];
    assign w_8_36 = data_operandA[28] & data_operandB[8];
    assign w_8_37 = data_operandA[29] & data_operandB[8];
    assign w_8_38 = data_operandA[30] & data_operandB[8];
    assign w_8_39 = ~(data_operandA[31] & data_operandB[8]);
    full_adder adder_8_8(.S(s_8_8), .Cout(c_8_8), .A(s_7_8), .B(w_8_8), .Cin(1'b0));
    full_adder adder_8_9(.S(s_8_9), .Cout(c_8_9), .A(s_7_9), .B(w_8_9), .Cin(c_8_8));
    full_adder adder_8_10(.S(s_8_10), .Cout(c_8_10), .A(s_7_10), .B(w_8_10), .Cin(c_8_9));
    full_adder adder_8_11(.S(s_8_11), .Cout(c_8_11), .A(s_7_11), .B(w_8_11), .Cin(c_8_10));
    full_adder adder_8_12(.S(s_8_12), .Cout(c_8_12), .A(s_7_12), .B(w_8_12), .Cin(c_8_11));
    full_adder adder_8_13(.S(s_8_13), .Cout(c_8_13), .A(s_7_13), .B(w_8_13), .Cin(c_8_12));
    full_adder adder_8_14(.S(s_8_14), .Cout(c_8_14), .A(s_7_14), .B(w_8_14), .Cin(c_8_13));
    full_adder adder_8_15(.S(s_8_15), .Cout(c_8_15), .A(s_7_15), .B(w_8_15), .Cin(c_8_14));
    full_adder adder_8_16(.S(s_8_16), .Cout(c_8_16), .A(s_7_16), .B(w_8_16), .Cin(c_8_15));
    full_adder adder_8_17(.S(s_8_17), .Cout(c_8_17), .A(s_7_17), .B(w_8_17), .Cin(c_8_16));
    full_adder adder_8_18(.S(s_8_18), .Cout(c_8_18), .A(s_7_18), .B(w_8_18), .Cin(c_8_17));
    full_adder adder_8_19(.S(s_8_19), .Cout(c_8_19), .A(s_7_19), .B(w_8_19), .Cin(c_8_18));
    full_adder adder_8_20(.S(s_8_20), .Cout(c_8_20), .A(s_7_20), .B(w_8_20), .Cin(c_8_19));
    full_adder adder_8_21(.S(s_8_21), .Cout(c_8_21), .A(s_7_21), .B(w_8_21), .Cin(c_8_20));
    full_adder adder_8_22(.S(s_8_22), .Cout(c_8_22), .A(s_7_22), .B(w_8_22), .Cin(c_8_21));
    full_adder adder_8_23(.S(s_8_23), .Cout(c_8_23), .A(s_7_23), .B(w_8_23), .Cin(c_8_22));
    full_adder adder_8_24(.S(s_8_24), .Cout(c_8_24), .A(s_7_24), .B(w_8_24), .Cin(c_8_23));
    full_adder adder_8_25(.S(s_8_25), .Cout(c_8_25), .A(s_7_25), .B(w_8_25), .Cin(c_8_24));
    full_adder adder_8_26(.S(s_8_26), .Cout(c_8_26), .A(s_7_26), .B(w_8_26), .Cin(c_8_25));
    full_adder adder_8_27(.S(s_8_27), .Cout(c_8_27), .A(s_7_27), .B(w_8_27), .Cin(c_8_26));
    full_adder adder_8_28(.S(s_8_28), .Cout(c_8_28), .A(s_7_28), .B(w_8_28), .Cin(c_8_27));
    full_adder adder_8_29(.S(s_8_29), .Cout(c_8_29), .A(s_7_29), .B(w_8_29), .Cin(c_8_28));
    full_adder adder_8_30(.S(s_8_30), .Cout(c_8_30), .A(s_7_30), .B(w_8_30), .Cin(c_8_29));
    full_adder adder_8_31(.S(s_8_31), .Cout(c_8_31), .A(s_7_31), .B(w_8_31), .Cin(c_8_30));
    full_adder adder_8_32(.S(s_8_32), .Cout(c_8_32), .A(s_7_32), .B(w_8_32), .Cin(c_8_31));
    full_adder adder_8_33(.S(s_8_33), .Cout(c_8_33), .A(s_7_33), .B(w_8_33), .Cin(c_8_32));
    full_adder adder_8_34(.S(s_8_34), .Cout(c_8_34), .A(s_7_34), .B(w_8_34), .Cin(c_8_33));
    full_adder adder_8_35(.S(s_8_35), .Cout(c_8_35), .A(s_7_35), .B(w_8_35), .Cin(c_8_34));
    full_adder adder_8_36(.S(s_8_36), .Cout(c_8_36), .A(s_7_36), .B(w_8_36), .Cin(c_8_35));
    full_adder adder_8_37(.S(s_8_37), .Cout(c_8_37), .A(s_7_37), .B(w_8_37), .Cin(c_8_36));
    full_adder adder_8_38(.S(s_8_38), .Cout(c_8_38), .A(s_7_38), .B(w_8_38), .Cin(c_8_37));
    full_adder adder_8_39(.S(s_8_39), .Cout(c_8_39), .A(c_7_38), .B(w_8_39), .Cin(c_8_38));
    assign result[8] = s_8_8;
    wire w_9_9, w_9_10, w_9_11, w_9_12, w_9_13, w_9_14, w_9_15, w_9_16, w_9_17, w_9_18, w_9_19, w_9_20, w_9_21, w_9_22, w_9_23, w_9_24, w_9_25, w_9_26, w_9_27, w_9_28, w_9_29, w_9_30, w_9_31, w_9_32, w_9_33, w_9_34, w_9_35, w_9_36, w_9_37, w_9_38, w_9_39, w_9_40;
    wire s_9_9, s_9_10, s_9_11, s_9_12, s_9_13, s_9_14, s_9_15, s_9_16, s_9_17, s_9_18, s_9_19, s_9_20, s_9_21, s_9_22, s_9_23, s_9_24, s_9_25, s_9_26, s_9_27, s_9_28, s_9_29, s_9_30, s_9_31, s_9_32, s_9_33, s_9_34, s_9_35, s_9_36, s_9_37, s_9_38, s_9_39, s_9_40;
    wire c_9_9, c_9_10, c_9_11, c_9_12, c_9_13, c_9_14, c_9_15, c_9_16, c_9_17, c_9_18, c_9_19, c_9_20, c_9_21, c_9_22, c_9_23, c_9_24, c_9_25, c_9_26, c_9_27, c_9_28, c_9_29, c_9_30, c_9_31, c_9_32, c_9_33, c_9_34, c_9_35, c_9_36, c_9_37, c_9_38, c_9_39, c_9_40;
    assign w_9_9 = data_operandA[0] & data_operandB[9];
    assign w_9_10 = data_operandA[1] & data_operandB[9];
    assign w_9_11 = data_operandA[2] & data_operandB[9];
    assign w_9_12 = data_operandA[3] & data_operandB[9];
    assign w_9_13 = data_operandA[4] & data_operandB[9];
    assign w_9_14 = data_operandA[5] & data_operandB[9];
    assign w_9_15 = data_operandA[6] & data_operandB[9];
    assign w_9_16 = data_operandA[7] & data_operandB[9];
    assign w_9_17 = data_operandA[8] & data_operandB[9];
    assign w_9_18 = data_operandA[9] & data_operandB[9];
    assign w_9_19 = data_operandA[10] & data_operandB[9];
    assign w_9_20 = data_operandA[11] & data_operandB[9];
    assign w_9_21 = data_operandA[12] & data_operandB[9];
    assign w_9_22 = data_operandA[13] & data_operandB[9];
    assign w_9_23 = data_operandA[14] & data_operandB[9];
    assign w_9_24 = data_operandA[15] & data_operandB[9];
    assign w_9_25 = data_operandA[16] & data_operandB[9];
    assign w_9_26 = data_operandA[17] & data_operandB[9];
    assign w_9_27 = data_operandA[18] & data_operandB[9];
    assign w_9_28 = data_operandA[19] & data_operandB[9];
    assign w_9_29 = data_operandA[20] & data_operandB[9];
    assign w_9_30 = data_operandA[21] & data_operandB[9];
    assign w_9_31 = data_operandA[22] & data_operandB[9];
    assign w_9_32 = data_operandA[23] & data_operandB[9];
    assign w_9_33 = data_operandA[24] & data_operandB[9];
    assign w_9_34 = data_operandA[25] & data_operandB[9];
    assign w_9_35 = data_operandA[26] & data_operandB[9];
    assign w_9_36 = data_operandA[27] & data_operandB[9];
    assign w_9_37 = data_operandA[28] & data_operandB[9];
    assign w_9_38 = data_operandA[29] & data_operandB[9];
    assign w_9_39 = data_operandA[30] & data_operandB[9];
    assign w_9_40 = ~(data_operandA[31] & data_operandB[9]);
    full_adder adder_9_9(.S(s_9_9), .Cout(c_9_9), .A(s_8_9), .B(w_9_9), .Cin(1'b0));
    full_adder adder_9_10(.S(s_9_10), .Cout(c_9_10), .A(s_8_10), .B(w_9_10), .Cin(c_9_9));
    full_adder adder_9_11(.S(s_9_11), .Cout(c_9_11), .A(s_8_11), .B(w_9_11), .Cin(c_9_10));
    full_adder adder_9_12(.S(s_9_12), .Cout(c_9_12), .A(s_8_12), .B(w_9_12), .Cin(c_9_11));
    full_adder adder_9_13(.S(s_9_13), .Cout(c_9_13), .A(s_8_13), .B(w_9_13), .Cin(c_9_12));
    full_adder adder_9_14(.S(s_9_14), .Cout(c_9_14), .A(s_8_14), .B(w_9_14), .Cin(c_9_13));
    full_adder adder_9_15(.S(s_9_15), .Cout(c_9_15), .A(s_8_15), .B(w_9_15), .Cin(c_9_14));
    full_adder adder_9_16(.S(s_9_16), .Cout(c_9_16), .A(s_8_16), .B(w_9_16), .Cin(c_9_15));
    full_adder adder_9_17(.S(s_9_17), .Cout(c_9_17), .A(s_8_17), .B(w_9_17), .Cin(c_9_16));
    full_adder adder_9_18(.S(s_9_18), .Cout(c_9_18), .A(s_8_18), .B(w_9_18), .Cin(c_9_17));
    full_adder adder_9_19(.S(s_9_19), .Cout(c_9_19), .A(s_8_19), .B(w_9_19), .Cin(c_9_18));
    full_adder adder_9_20(.S(s_9_20), .Cout(c_9_20), .A(s_8_20), .B(w_9_20), .Cin(c_9_19));
    full_adder adder_9_21(.S(s_9_21), .Cout(c_9_21), .A(s_8_21), .B(w_9_21), .Cin(c_9_20));
    full_adder adder_9_22(.S(s_9_22), .Cout(c_9_22), .A(s_8_22), .B(w_9_22), .Cin(c_9_21));
    full_adder adder_9_23(.S(s_9_23), .Cout(c_9_23), .A(s_8_23), .B(w_9_23), .Cin(c_9_22));
    full_adder adder_9_24(.S(s_9_24), .Cout(c_9_24), .A(s_8_24), .B(w_9_24), .Cin(c_9_23));
    full_adder adder_9_25(.S(s_9_25), .Cout(c_9_25), .A(s_8_25), .B(w_9_25), .Cin(c_9_24));
    full_adder adder_9_26(.S(s_9_26), .Cout(c_9_26), .A(s_8_26), .B(w_9_26), .Cin(c_9_25));
    full_adder adder_9_27(.S(s_9_27), .Cout(c_9_27), .A(s_8_27), .B(w_9_27), .Cin(c_9_26));
    full_adder adder_9_28(.S(s_9_28), .Cout(c_9_28), .A(s_8_28), .B(w_9_28), .Cin(c_9_27));
    full_adder adder_9_29(.S(s_9_29), .Cout(c_9_29), .A(s_8_29), .B(w_9_29), .Cin(c_9_28));
    full_adder adder_9_30(.S(s_9_30), .Cout(c_9_30), .A(s_8_30), .B(w_9_30), .Cin(c_9_29));
    full_adder adder_9_31(.S(s_9_31), .Cout(c_9_31), .A(s_8_31), .B(w_9_31), .Cin(c_9_30));
    full_adder adder_9_32(.S(s_9_32), .Cout(c_9_32), .A(s_8_32), .B(w_9_32), .Cin(c_9_31));
    full_adder adder_9_33(.S(s_9_33), .Cout(c_9_33), .A(s_8_33), .B(w_9_33), .Cin(c_9_32));
    full_adder adder_9_34(.S(s_9_34), .Cout(c_9_34), .A(s_8_34), .B(w_9_34), .Cin(c_9_33));
    full_adder adder_9_35(.S(s_9_35), .Cout(c_9_35), .A(s_8_35), .B(w_9_35), .Cin(c_9_34));
    full_adder adder_9_36(.S(s_9_36), .Cout(c_9_36), .A(s_8_36), .B(w_9_36), .Cin(c_9_35));
    full_adder adder_9_37(.S(s_9_37), .Cout(c_9_37), .A(s_8_37), .B(w_9_37), .Cin(c_9_36));
    full_adder adder_9_38(.S(s_9_38), .Cout(c_9_38), .A(s_8_38), .B(w_9_38), .Cin(c_9_37));
    full_adder adder_9_39(.S(s_9_39), .Cout(c_9_39), .A(s_8_39), .B(w_9_39), .Cin(c_9_38));
    full_adder adder_9_40(.S(s_9_40), .Cout(c_9_40), .A(c_8_39), .B(w_9_40), .Cin(c_9_39));
    assign result[9] = s_9_9;
    wire w_10_10, w_10_11, w_10_12, w_10_13, w_10_14, w_10_15, w_10_16, w_10_17, w_10_18, w_10_19, w_10_20, w_10_21, w_10_22, w_10_23, w_10_24, w_10_25, w_10_26, w_10_27, w_10_28, w_10_29, w_10_30, w_10_31, w_10_32, w_10_33, w_10_34, w_10_35, w_10_36, w_10_37, w_10_38, w_10_39, w_10_40, w_10_41;
    wire s_10_10, s_10_11, s_10_12, s_10_13, s_10_14, s_10_15, s_10_16, s_10_17, s_10_18, s_10_19, s_10_20, s_10_21, s_10_22, s_10_23, s_10_24, s_10_25, s_10_26, s_10_27, s_10_28, s_10_29, s_10_30, s_10_31, s_10_32, s_10_33, s_10_34, s_10_35, s_10_36, s_10_37, s_10_38, s_10_39, s_10_40, s_10_41;
    wire c_10_10, c_10_11, c_10_12, c_10_13, c_10_14, c_10_15, c_10_16, c_10_17, c_10_18, c_10_19, c_10_20, c_10_21, c_10_22, c_10_23, c_10_24, c_10_25, c_10_26, c_10_27, c_10_28, c_10_29, c_10_30, c_10_31, c_10_32, c_10_33, c_10_34, c_10_35, c_10_36, c_10_37, c_10_38, c_10_39, c_10_40, c_10_41;
    assign w_10_10 = data_operandA[0] & data_operandB[10];
    assign w_10_11 = data_operandA[1] & data_operandB[10];
    assign w_10_12 = data_operandA[2] & data_operandB[10];
    assign w_10_13 = data_operandA[3] & data_operandB[10];
    assign w_10_14 = data_operandA[4] & data_operandB[10];
    assign w_10_15 = data_operandA[5] & data_operandB[10];
    assign w_10_16 = data_operandA[6] & data_operandB[10];
    assign w_10_17 = data_operandA[7] & data_operandB[10];
    assign w_10_18 = data_operandA[8] & data_operandB[10];
    assign w_10_19 = data_operandA[9] & data_operandB[10];
    assign w_10_20 = data_operandA[10] & data_operandB[10];
    assign w_10_21 = data_operandA[11] & data_operandB[10];
    assign w_10_22 = data_operandA[12] & data_operandB[10];
    assign w_10_23 = data_operandA[13] & data_operandB[10];
    assign w_10_24 = data_operandA[14] & data_operandB[10];
    assign w_10_25 = data_operandA[15] & data_operandB[10];
    assign w_10_26 = data_operandA[16] & data_operandB[10];
    assign w_10_27 = data_operandA[17] & data_operandB[10];
    assign w_10_28 = data_operandA[18] & data_operandB[10];
    assign w_10_29 = data_operandA[19] & data_operandB[10];
    assign w_10_30 = data_operandA[20] & data_operandB[10];
    assign w_10_31 = data_operandA[21] & data_operandB[10];
    assign w_10_32 = data_operandA[22] & data_operandB[10];
    assign w_10_33 = data_operandA[23] & data_operandB[10];
    assign w_10_34 = data_operandA[24] & data_operandB[10];
    assign w_10_35 = data_operandA[25] & data_operandB[10];
    assign w_10_36 = data_operandA[26] & data_operandB[10];
    assign w_10_37 = data_operandA[27] & data_operandB[10];
    assign w_10_38 = data_operandA[28] & data_operandB[10];
    assign w_10_39 = data_operandA[29] & data_operandB[10];
    assign w_10_40 = data_operandA[30] & data_operandB[10];
    assign w_10_41 = ~(data_operandA[31] & data_operandB[10]);
    full_adder adder_10_10(.S(s_10_10), .Cout(c_10_10), .A(s_9_10), .B(w_10_10), .Cin(1'b0));
    full_adder adder_10_11(.S(s_10_11), .Cout(c_10_11), .A(s_9_11), .B(w_10_11), .Cin(c_10_10));
    full_adder adder_10_12(.S(s_10_12), .Cout(c_10_12), .A(s_9_12), .B(w_10_12), .Cin(c_10_11));
    full_adder adder_10_13(.S(s_10_13), .Cout(c_10_13), .A(s_9_13), .B(w_10_13), .Cin(c_10_12));
    full_adder adder_10_14(.S(s_10_14), .Cout(c_10_14), .A(s_9_14), .B(w_10_14), .Cin(c_10_13));
    full_adder adder_10_15(.S(s_10_15), .Cout(c_10_15), .A(s_9_15), .B(w_10_15), .Cin(c_10_14));
    full_adder adder_10_16(.S(s_10_16), .Cout(c_10_16), .A(s_9_16), .B(w_10_16), .Cin(c_10_15));
    full_adder adder_10_17(.S(s_10_17), .Cout(c_10_17), .A(s_9_17), .B(w_10_17), .Cin(c_10_16));
    full_adder adder_10_18(.S(s_10_18), .Cout(c_10_18), .A(s_9_18), .B(w_10_18), .Cin(c_10_17));
    full_adder adder_10_19(.S(s_10_19), .Cout(c_10_19), .A(s_9_19), .B(w_10_19), .Cin(c_10_18));
    full_adder adder_10_20(.S(s_10_20), .Cout(c_10_20), .A(s_9_20), .B(w_10_20), .Cin(c_10_19));
    full_adder adder_10_21(.S(s_10_21), .Cout(c_10_21), .A(s_9_21), .B(w_10_21), .Cin(c_10_20));
    full_adder adder_10_22(.S(s_10_22), .Cout(c_10_22), .A(s_9_22), .B(w_10_22), .Cin(c_10_21));
    full_adder adder_10_23(.S(s_10_23), .Cout(c_10_23), .A(s_9_23), .B(w_10_23), .Cin(c_10_22));
    full_adder adder_10_24(.S(s_10_24), .Cout(c_10_24), .A(s_9_24), .B(w_10_24), .Cin(c_10_23));
    full_adder adder_10_25(.S(s_10_25), .Cout(c_10_25), .A(s_9_25), .B(w_10_25), .Cin(c_10_24));
    full_adder adder_10_26(.S(s_10_26), .Cout(c_10_26), .A(s_9_26), .B(w_10_26), .Cin(c_10_25));
    full_adder adder_10_27(.S(s_10_27), .Cout(c_10_27), .A(s_9_27), .B(w_10_27), .Cin(c_10_26));
    full_adder adder_10_28(.S(s_10_28), .Cout(c_10_28), .A(s_9_28), .B(w_10_28), .Cin(c_10_27));
    full_adder adder_10_29(.S(s_10_29), .Cout(c_10_29), .A(s_9_29), .B(w_10_29), .Cin(c_10_28));
    full_adder adder_10_30(.S(s_10_30), .Cout(c_10_30), .A(s_9_30), .B(w_10_30), .Cin(c_10_29));
    full_adder adder_10_31(.S(s_10_31), .Cout(c_10_31), .A(s_9_31), .B(w_10_31), .Cin(c_10_30));
    full_adder adder_10_32(.S(s_10_32), .Cout(c_10_32), .A(s_9_32), .B(w_10_32), .Cin(c_10_31));
    full_adder adder_10_33(.S(s_10_33), .Cout(c_10_33), .A(s_9_33), .B(w_10_33), .Cin(c_10_32));
    full_adder adder_10_34(.S(s_10_34), .Cout(c_10_34), .A(s_9_34), .B(w_10_34), .Cin(c_10_33));
    full_adder adder_10_35(.S(s_10_35), .Cout(c_10_35), .A(s_9_35), .B(w_10_35), .Cin(c_10_34));
    full_adder adder_10_36(.S(s_10_36), .Cout(c_10_36), .A(s_9_36), .B(w_10_36), .Cin(c_10_35));
    full_adder adder_10_37(.S(s_10_37), .Cout(c_10_37), .A(s_9_37), .B(w_10_37), .Cin(c_10_36));
    full_adder adder_10_38(.S(s_10_38), .Cout(c_10_38), .A(s_9_38), .B(w_10_38), .Cin(c_10_37));
    full_adder adder_10_39(.S(s_10_39), .Cout(c_10_39), .A(s_9_39), .B(w_10_39), .Cin(c_10_38));
    full_adder adder_10_40(.S(s_10_40), .Cout(c_10_40), .A(s_9_40), .B(w_10_40), .Cin(c_10_39));
    full_adder adder_10_41(.S(s_10_41), .Cout(c_10_41), .A(c_9_40), .B(w_10_41), .Cin(c_10_40));
    assign result[10] = s_10_10;
    wire w_11_11, w_11_12, w_11_13, w_11_14, w_11_15, w_11_16, w_11_17, w_11_18, w_11_19, w_11_20, w_11_21, w_11_22, w_11_23, w_11_24, w_11_25, w_11_26, w_11_27, w_11_28, w_11_29, w_11_30, w_11_31, w_11_32, w_11_33, w_11_34, w_11_35, w_11_36, w_11_37, w_11_38, w_11_39, w_11_40, w_11_41, w_11_42;
    wire s_11_11, s_11_12, s_11_13, s_11_14, s_11_15, s_11_16, s_11_17, s_11_18, s_11_19, s_11_20, s_11_21, s_11_22, s_11_23, s_11_24, s_11_25, s_11_26, s_11_27, s_11_28, s_11_29, s_11_30, s_11_31, s_11_32, s_11_33, s_11_34, s_11_35, s_11_36, s_11_37, s_11_38, s_11_39, s_11_40, s_11_41, s_11_42;
    wire c_11_11, c_11_12, c_11_13, c_11_14, c_11_15, c_11_16, c_11_17, c_11_18, c_11_19, c_11_20, c_11_21, c_11_22, c_11_23, c_11_24, c_11_25, c_11_26, c_11_27, c_11_28, c_11_29, c_11_30, c_11_31, c_11_32, c_11_33, c_11_34, c_11_35, c_11_36, c_11_37, c_11_38, c_11_39, c_11_40, c_11_41, c_11_42;
    assign w_11_11 = data_operandA[0] & data_operandB[11];
    assign w_11_12 = data_operandA[1] & data_operandB[11];
    assign w_11_13 = data_operandA[2] & data_operandB[11];
    assign w_11_14 = data_operandA[3] & data_operandB[11];
    assign w_11_15 = data_operandA[4] & data_operandB[11];
    assign w_11_16 = data_operandA[5] & data_operandB[11];
    assign w_11_17 = data_operandA[6] & data_operandB[11];
    assign w_11_18 = data_operandA[7] & data_operandB[11];
    assign w_11_19 = data_operandA[8] & data_operandB[11];
    assign w_11_20 = data_operandA[9] & data_operandB[11];
    assign w_11_21 = data_operandA[10] & data_operandB[11];
    assign w_11_22 = data_operandA[11] & data_operandB[11];
    assign w_11_23 = data_operandA[12] & data_operandB[11];
    assign w_11_24 = data_operandA[13] & data_operandB[11];
    assign w_11_25 = data_operandA[14] & data_operandB[11];
    assign w_11_26 = data_operandA[15] & data_operandB[11];
    assign w_11_27 = data_operandA[16] & data_operandB[11];
    assign w_11_28 = data_operandA[17] & data_operandB[11];
    assign w_11_29 = data_operandA[18] & data_operandB[11];
    assign w_11_30 = data_operandA[19] & data_operandB[11];
    assign w_11_31 = data_operandA[20] & data_operandB[11];
    assign w_11_32 = data_operandA[21] & data_operandB[11];
    assign w_11_33 = data_operandA[22] & data_operandB[11];
    assign w_11_34 = data_operandA[23] & data_operandB[11];
    assign w_11_35 = data_operandA[24] & data_operandB[11];
    assign w_11_36 = data_operandA[25] & data_operandB[11];
    assign w_11_37 = data_operandA[26] & data_operandB[11];
    assign w_11_38 = data_operandA[27] & data_operandB[11];
    assign w_11_39 = data_operandA[28] & data_operandB[11];
    assign w_11_40 = data_operandA[29] & data_operandB[11];
    assign w_11_41 = data_operandA[30] & data_operandB[11];
    assign w_11_42 = ~(data_operandA[31] & data_operandB[11]);
    full_adder adder_11_11(.S(s_11_11), .Cout(c_11_11), .A(s_10_11), .B(w_11_11), .Cin(1'b0));
    full_adder adder_11_12(.S(s_11_12), .Cout(c_11_12), .A(s_10_12), .B(w_11_12), .Cin(c_11_11));
    full_adder adder_11_13(.S(s_11_13), .Cout(c_11_13), .A(s_10_13), .B(w_11_13), .Cin(c_11_12));
    full_adder adder_11_14(.S(s_11_14), .Cout(c_11_14), .A(s_10_14), .B(w_11_14), .Cin(c_11_13));
    full_adder adder_11_15(.S(s_11_15), .Cout(c_11_15), .A(s_10_15), .B(w_11_15), .Cin(c_11_14));
    full_adder adder_11_16(.S(s_11_16), .Cout(c_11_16), .A(s_10_16), .B(w_11_16), .Cin(c_11_15));
    full_adder adder_11_17(.S(s_11_17), .Cout(c_11_17), .A(s_10_17), .B(w_11_17), .Cin(c_11_16));
    full_adder adder_11_18(.S(s_11_18), .Cout(c_11_18), .A(s_10_18), .B(w_11_18), .Cin(c_11_17));
    full_adder adder_11_19(.S(s_11_19), .Cout(c_11_19), .A(s_10_19), .B(w_11_19), .Cin(c_11_18));
    full_adder adder_11_20(.S(s_11_20), .Cout(c_11_20), .A(s_10_20), .B(w_11_20), .Cin(c_11_19));
    full_adder adder_11_21(.S(s_11_21), .Cout(c_11_21), .A(s_10_21), .B(w_11_21), .Cin(c_11_20));
    full_adder adder_11_22(.S(s_11_22), .Cout(c_11_22), .A(s_10_22), .B(w_11_22), .Cin(c_11_21));
    full_adder adder_11_23(.S(s_11_23), .Cout(c_11_23), .A(s_10_23), .B(w_11_23), .Cin(c_11_22));
    full_adder adder_11_24(.S(s_11_24), .Cout(c_11_24), .A(s_10_24), .B(w_11_24), .Cin(c_11_23));
    full_adder adder_11_25(.S(s_11_25), .Cout(c_11_25), .A(s_10_25), .B(w_11_25), .Cin(c_11_24));
    full_adder adder_11_26(.S(s_11_26), .Cout(c_11_26), .A(s_10_26), .B(w_11_26), .Cin(c_11_25));
    full_adder adder_11_27(.S(s_11_27), .Cout(c_11_27), .A(s_10_27), .B(w_11_27), .Cin(c_11_26));
    full_adder adder_11_28(.S(s_11_28), .Cout(c_11_28), .A(s_10_28), .B(w_11_28), .Cin(c_11_27));
    full_adder adder_11_29(.S(s_11_29), .Cout(c_11_29), .A(s_10_29), .B(w_11_29), .Cin(c_11_28));
    full_adder adder_11_30(.S(s_11_30), .Cout(c_11_30), .A(s_10_30), .B(w_11_30), .Cin(c_11_29));
    full_adder adder_11_31(.S(s_11_31), .Cout(c_11_31), .A(s_10_31), .B(w_11_31), .Cin(c_11_30));
    full_adder adder_11_32(.S(s_11_32), .Cout(c_11_32), .A(s_10_32), .B(w_11_32), .Cin(c_11_31));
    full_adder adder_11_33(.S(s_11_33), .Cout(c_11_33), .A(s_10_33), .B(w_11_33), .Cin(c_11_32));
    full_adder adder_11_34(.S(s_11_34), .Cout(c_11_34), .A(s_10_34), .B(w_11_34), .Cin(c_11_33));
    full_adder adder_11_35(.S(s_11_35), .Cout(c_11_35), .A(s_10_35), .B(w_11_35), .Cin(c_11_34));
    full_adder adder_11_36(.S(s_11_36), .Cout(c_11_36), .A(s_10_36), .B(w_11_36), .Cin(c_11_35));
    full_adder adder_11_37(.S(s_11_37), .Cout(c_11_37), .A(s_10_37), .B(w_11_37), .Cin(c_11_36));
    full_adder adder_11_38(.S(s_11_38), .Cout(c_11_38), .A(s_10_38), .B(w_11_38), .Cin(c_11_37));
    full_adder adder_11_39(.S(s_11_39), .Cout(c_11_39), .A(s_10_39), .B(w_11_39), .Cin(c_11_38));
    full_adder adder_11_40(.S(s_11_40), .Cout(c_11_40), .A(s_10_40), .B(w_11_40), .Cin(c_11_39));
    full_adder adder_11_41(.S(s_11_41), .Cout(c_11_41), .A(s_10_41), .B(w_11_41), .Cin(c_11_40));
    full_adder adder_11_42(.S(s_11_42), .Cout(c_11_42), .A(c_10_41), .B(w_11_42), .Cin(c_11_41));
    assign result[11] = s_11_11;
    wire w_12_12, w_12_13, w_12_14, w_12_15, w_12_16, w_12_17, w_12_18, w_12_19, w_12_20, w_12_21, w_12_22, w_12_23, w_12_24, w_12_25, w_12_26, w_12_27, w_12_28, w_12_29, w_12_30, w_12_31, w_12_32, w_12_33, w_12_34, w_12_35, w_12_36, w_12_37, w_12_38, w_12_39, w_12_40, w_12_41, w_12_42, w_12_43;
    wire s_12_12, s_12_13, s_12_14, s_12_15, s_12_16, s_12_17, s_12_18, s_12_19, s_12_20, s_12_21, s_12_22, s_12_23, s_12_24, s_12_25, s_12_26, s_12_27, s_12_28, s_12_29, s_12_30, s_12_31, s_12_32, s_12_33, s_12_34, s_12_35, s_12_36, s_12_37, s_12_38, s_12_39, s_12_40, s_12_41, s_12_42, s_12_43;
    wire c_12_12, c_12_13, c_12_14, c_12_15, c_12_16, c_12_17, c_12_18, c_12_19, c_12_20, c_12_21, c_12_22, c_12_23, c_12_24, c_12_25, c_12_26, c_12_27, c_12_28, c_12_29, c_12_30, c_12_31, c_12_32, c_12_33, c_12_34, c_12_35, c_12_36, c_12_37, c_12_38, c_12_39, c_12_40, c_12_41, c_12_42, c_12_43;
    assign w_12_12 = data_operandA[0] & data_operandB[12];
    assign w_12_13 = data_operandA[1] & data_operandB[12];
    assign w_12_14 = data_operandA[2] & data_operandB[12];
    assign w_12_15 = data_operandA[3] & data_operandB[12];
    assign w_12_16 = data_operandA[4] & data_operandB[12];
    assign w_12_17 = data_operandA[5] & data_operandB[12];
    assign w_12_18 = data_operandA[6] & data_operandB[12];
    assign w_12_19 = data_operandA[7] & data_operandB[12];
    assign w_12_20 = data_operandA[8] & data_operandB[12];
    assign w_12_21 = data_operandA[9] & data_operandB[12];
    assign w_12_22 = data_operandA[10] & data_operandB[12];
    assign w_12_23 = data_operandA[11] & data_operandB[12];
    assign w_12_24 = data_operandA[12] & data_operandB[12];
    assign w_12_25 = data_operandA[13] & data_operandB[12];
    assign w_12_26 = data_operandA[14] & data_operandB[12];
    assign w_12_27 = data_operandA[15] & data_operandB[12];
    assign w_12_28 = data_operandA[16] & data_operandB[12];
    assign w_12_29 = data_operandA[17] & data_operandB[12];
    assign w_12_30 = data_operandA[18] & data_operandB[12];
    assign w_12_31 = data_operandA[19] & data_operandB[12];
    assign w_12_32 = data_operandA[20] & data_operandB[12];
    assign w_12_33 = data_operandA[21] & data_operandB[12];
    assign w_12_34 = data_operandA[22] & data_operandB[12];
    assign w_12_35 = data_operandA[23] & data_operandB[12];
    assign w_12_36 = data_operandA[24] & data_operandB[12];
    assign w_12_37 = data_operandA[25] & data_operandB[12];
    assign w_12_38 = data_operandA[26] & data_operandB[12];
    assign w_12_39 = data_operandA[27] & data_operandB[12];
    assign w_12_40 = data_operandA[28] & data_operandB[12];
    assign w_12_41 = data_operandA[29] & data_operandB[12];
    assign w_12_42 = data_operandA[30] & data_operandB[12];
    assign w_12_43 = ~(data_operandA[31] & data_operandB[12]);
    full_adder adder_12_12(.S(s_12_12), .Cout(c_12_12), .A(s_11_12), .B(w_12_12), .Cin(1'b0));
    full_adder adder_12_13(.S(s_12_13), .Cout(c_12_13), .A(s_11_13), .B(w_12_13), .Cin(c_12_12));
    full_adder adder_12_14(.S(s_12_14), .Cout(c_12_14), .A(s_11_14), .B(w_12_14), .Cin(c_12_13));
    full_adder adder_12_15(.S(s_12_15), .Cout(c_12_15), .A(s_11_15), .B(w_12_15), .Cin(c_12_14));
    full_adder adder_12_16(.S(s_12_16), .Cout(c_12_16), .A(s_11_16), .B(w_12_16), .Cin(c_12_15));
    full_adder adder_12_17(.S(s_12_17), .Cout(c_12_17), .A(s_11_17), .B(w_12_17), .Cin(c_12_16));
    full_adder adder_12_18(.S(s_12_18), .Cout(c_12_18), .A(s_11_18), .B(w_12_18), .Cin(c_12_17));
    full_adder adder_12_19(.S(s_12_19), .Cout(c_12_19), .A(s_11_19), .B(w_12_19), .Cin(c_12_18));
    full_adder adder_12_20(.S(s_12_20), .Cout(c_12_20), .A(s_11_20), .B(w_12_20), .Cin(c_12_19));
    full_adder adder_12_21(.S(s_12_21), .Cout(c_12_21), .A(s_11_21), .B(w_12_21), .Cin(c_12_20));
    full_adder adder_12_22(.S(s_12_22), .Cout(c_12_22), .A(s_11_22), .B(w_12_22), .Cin(c_12_21));
    full_adder adder_12_23(.S(s_12_23), .Cout(c_12_23), .A(s_11_23), .B(w_12_23), .Cin(c_12_22));
    full_adder adder_12_24(.S(s_12_24), .Cout(c_12_24), .A(s_11_24), .B(w_12_24), .Cin(c_12_23));
    full_adder adder_12_25(.S(s_12_25), .Cout(c_12_25), .A(s_11_25), .B(w_12_25), .Cin(c_12_24));
    full_adder adder_12_26(.S(s_12_26), .Cout(c_12_26), .A(s_11_26), .B(w_12_26), .Cin(c_12_25));
    full_adder adder_12_27(.S(s_12_27), .Cout(c_12_27), .A(s_11_27), .B(w_12_27), .Cin(c_12_26));
    full_adder adder_12_28(.S(s_12_28), .Cout(c_12_28), .A(s_11_28), .B(w_12_28), .Cin(c_12_27));
    full_adder adder_12_29(.S(s_12_29), .Cout(c_12_29), .A(s_11_29), .B(w_12_29), .Cin(c_12_28));
    full_adder adder_12_30(.S(s_12_30), .Cout(c_12_30), .A(s_11_30), .B(w_12_30), .Cin(c_12_29));
    full_adder adder_12_31(.S(s_12_31), .Cout(c_12_31), .A(s_11_31), .B(w_12_31), .Cin(c_12_30));
    full_adder adder_12_32(.S(s_12_32), .Cout(c_12_32), .A(s_11_32), .B(w_12_32), .Cin(c_12_31));
    full_adder adder_12_33(.S(s_12_33), .Cout(c_12_33), .A(s_11_33), .B(w_12_33), .Cin(c_12_32));
    full_adder adder_12_34(.S(s_12_34), .Cout(c_12_34), .A(s_11_34), .B(w_12_34), .Cin(c_12_33));
    full_adder adder_12_35(.S(s_12_35), .Cout(c_12_35), .A(s_11_35), .B(w_12_35), .Cin(c_12_34));
    full_adder adder_12_36(.S(s_12_36), .Cout(c_12_36), .A(s_11_36), .B(w_12_36), .Cin(c_12_35));
    full_adder adder_12_37(.S(s_12_37), .Cout(c_12_37), .A(s_11_37), .B(w_12_37), .Cin(c_12_36));
    full_adder adder_12_38(.S(s_12_38), .Cout(c_12_38), .A(s_11_38), .B(w_12_38), .Cin(c_12_37));
    full_adder adder_12_39(.S(s_12_39), .Cout(c_12_39), .A(s_11_39), .B(w_12_39), .Cin(c_12_38));
    full_adder adder_12_40(.S(s_12_40), .Cout(c_12_40), .A(s_11_40), .B(w_12_40), .Cin(c_12_39));
    full_adder adder_12_41(.S(s_12_41), .Cout(c_12_41), .A(s_11_41), .B(w_12_41), .Cin(c_12_40));
    full_adder adder_12_42(.S(s_12_42), .Cout(c_12_42), .A(s_11_42), .B(w_12_42), .Cin(c_12_41));
    full_adder adder_12_43(.S(s_12_43), .Cout(c_12_43), .A(c_11_42), .B(w_12_43), .Cin(c_12_42));
    assign result[12] = s_12_12;
    wire w_13_13, w_13_14, w_13_15, w_13_16, w_13_17, w_13_18, w_13_19, w_13_20, w_13_21, w_13_22, w_13_23, w_13_24, w_13_25, w_13_26, w_13_27, w_13_28, w_13_29, w_13_30, w_13_31, w_13_32, w_13_33, w_13_34, w_13_35, w_13_36, w_13_37, w_13_38, w_13_39, w_13_40, w_13_41, w_13_42, w_13_43, w_13_44;
    wire s_13_13, s_13_14, s_13_15, s_13_16, s_13_17, s_13_18, s_13_19, s_13_20, s_13_21, s_13_22, s_13_23, s_13_24, s_13_25, s_13_26, s_13_27, s_13_28, s_13_29, s_13_30, s_13_31, s_13_32, s_13_33, s_13_34, s_13_35, s_13_36, s_13_37, s_13_38, s_13_39, s_13_40, s_13_41, s_13_42, s_13_43, s_13_44;
    wire c_13_13, c_13_14, c_13_15, c_13_16, c_13_17, c_13_18, c_13_19, c_13_20, c_13_21, c_13_22, c_13_23, c_13_24, c_13_25, c_13_26, c_13_27, c_13_28, c_13_29, c_13_30, c_13_31, c_13_32, c_13_33, c_13_34, c_13_35, c_13_36, c_13_37, c_13_38, c_13_39, c_13_40, c_13_41, c_13_42, c_13_43, c_13_44;
    assign w_13_13 = data_operandA[0] & data_operandB[13];
    assign w_13_14 = data_operandA[1] & data_operandB[13];
    assign w_13_15 = data_operandA[2] & data_operandB[13];
    assign w_13_16 = data_operandA[3] & data_operandB[13];
    assign w_13_17 = data_operandA[4] & data_operandB[13];
    assign w_13_18 = data_operandA[5] & data_operandB[13];
    assign w_13_19 = data_operandA[6] & data_operandB[13];
    assign w_13_20 = data_operandA[7] & data_operandB[13];
    assign w_13_21 = data_operandA[8] & data_operandB[13];
    assign w_13_22 = data_operandA[9] & data_operandB[13];
    assign w_13_23 = data_operandA[10] & data_operandB[13];
    assign w_13_24 = data_operandA[11] & data_operandB[13];
    assign w_13_25 = data_operandA[12] & data_operandB[13];
    assign w_13_26 = data_operandA[13] & data_operandB[13];
    assign w_13_27 = data_operandA[14] & data_operandB[13];
    assign w_13_28 = data_operandA[15] & data_operandB[13];
    assign w_13_29 = data_operandA[16] & data_operandB[13];
    assign w_13_30 = data_operandA[17] & data_operandB[13];
    assign w_13_31 = data_operandA[18] & data_operandB[13];
    assign w_13_32 = data_operandA[19] & data_operandB[13];
    assign w_13_33 = data_operandA[20] & data_operandB[13];
    assign w_13_34 = data_operandA[21] & data_operandB[13];
    assign w_13_35 = data_operandA[22] & data_operandB[13];
    assign w_13_36 = data_operandA[23] & data_operandB[13];
    assign w_13_37 = data_operandA[24] & data_operandB[13];
    assign w_13_38 = data_operandA[25] & data_operandB[13];
    assign w_13_39 = data_operandA[26] & data_operandB[13];
    assign w_13_40 = data_operandA[27] & data_operandB[13];
    assign w_13_41 = data_operandA[28] & data_operandB[13];
    assign w_13_42 = data_operandA[29] & data_operandB[13];
    assign w_13_43 = data_operandA[30] & data_operandB[13];
    assign w_13_44 = ~(data_operandA[31] & data_operandB[13]);
    full_adder adder_13_13(.S(s_13_13), .Cout(c_13_13), .A(s_12_13), .B(w_13_13), .Cin(1'b0));
    full_adder adder_13_14(.S(s_13_14), .Cout(c_13_14), .A(s_12_14), .B(w_13_14), .Cin(c_13_13));
    full_adder adder_13_15(.S(s_13_15), .Cout(c_13_15), .A(s_12_15), .B(w_13_15), .Cin(c_13_14));
    full_adder adder_13_16(.S(s_13_16), .Cout(c_13_16), .A(s_12_16), .B(w_13_16), .Cin(c_13_15));
    full_adder adder_13_17(.S(s_13_17), .Cout(c_13_17), .A(s_12_17), .B(w_13_17), .Cin(c_13_16));
    full_adder adder_13_18(.S(s_13_18), .Cout(c_13_18), .A(s_12_18), .B(w_13_18), .Cin(c_13_17));
    full_adder adder_13_19(.S(s_13_19), .Cout(c_13_19), .A(s_12_19), .B(w_13_19), .Cin(c_13_18));
    full_adder adder_13_20(.S(s_13_20), .Cout(c_13_20), .A(s_12_20), .B(w_13_20), .Cin(c_13_19));
    full_adder adder_13_21(.S(s_13_21), .Cout(c_13_21), .A(s_12_21), .B(w_13_21), .Cin(c_13_20));
    full_adder adder_13_22(.S(s_13_22), .Cout(c_13_22), .A(s_12_22), .B(w_13_22), .Cin(c_13_21));
    full_adder adder_13_23(.S(s_13_23), .Cout(c_13_23), .A(s_12_23), .B(w_13_23), .Cin(c_13_22));
    full_adder adder_13_24(.S(s_13_24), .Cout(c_13_24), .A(s_12_24), .B(w_13_24), .Cin(c_13_23));
    full_adder adder_13_25(.S(s_13_25), .Cout(c_13_25), .A(s_12_25), .B(w_13_25), .Cin(c_13_24));
    full_adder adder_13_26(.S(s_13_26), .Cout(c_13_26), .A(s_12_26), .B(w_13_26), .Cin(c_13_25));
    full_adder adder_13_27(.S(s_13_27), .Cout(c_13_27), .A(s_12_27), .B(w_13_27), .Cin(c_13_26));
    full_adder adder_13_28(.S(s_13_28), .Cout(c_13_28), .A(s_12_28), .B(w_13_28), .Cin(c_13_27));
    full_adder adder_13_29(.S(s_13_29), .Cout(c_13_29), .A(s_12_29), .B(w_13_29), .Cin(c_13_28));
    full_adder adder_13_30(.S(s_13_30), .Cout(c_13_30), .A(s_12_30), .B(w_13_30), .Cin(c_13_29));
    full_adder adder_13_31(.S(s_13_31), .Cout(c_13_31), .A(s_12_31), .B(w_13_31), .Cin(c_13_30));
    full_adder adder_13_32(.S(s_13_32), .Cout(c_13_32), .A(s_12_32), .B(w_13_32), .Cin(c_13_31));
    full_adder adder_13_33(.S(s_13_33), .Cout(c_13_33), .A(s_12_33), .B(w_13_33), .Cin(c_13_32));
    full_adder adder_13_34(.S(s_13_34), .Cout(c_13_34), .A(s_12_34), .B(w_13_34), .Cin(c_13_33));
    full_adder adder_13_35(.S(s_13_35), .Cout(c_13_35), .A(s_12_35), .B(w_13_35), .Cin(c_13_34));
    full_adder adder_13_36(.S(s_13_36), .Cout(c_13_36), .A(s_12_36), .B(w_13_36), .Cin(c_13_35));
    full_adder adder_13_37(.S(s_13_37), .Cout(c_13_37), .A(s_12_37), .B(w_13_37), .Cin(c_13_36));
    full_adder adder_13_38(.S(s_13_38), .Cout(c_13_38), .A(s_12_38), .B(w_13_38), .Cin(c_13_37));
    full_adder adder_13_39(.S(s_13_39), .Cout(c_13_39), .A(s_12_39), .B(w_13_39), .Cin(c_13_38));
    full_adder adder_13_40(.S(s_13_40), .Cout(c_13_40), .A(s_12_40), .B(w_13_40), .Cin(c_13_39));
    full_adder adder_13_41(.S(s_13_41), .Cout(c_13_41), .A(s_12_41), .B(w_13_41), .Cin(c_13_40));
    full_adder adder_13_42(.S(s_13_42), .Cout(c_13_42), .A(s_12_42), .B(w_13_42), .Cin(c_13_41));
    full_adder adder_13_43(.S(s_13_43), .Cout(c_13_43), .A(s_12_43), .B(w_13_43), .Cin(c_13_42));
    full_adder adder_13_44(.S(s_13_44), .Cout(c_13_44), .A(c_12_43), .B(w_13_44), .Cin(c_13_43));
    assign result[13] = s_13_13;
    wire w_14_14, w_14_15, w_14_16, w_14_17, w_14_18, w_14_19, w_14_20, w_14_21, w_14_22, w_14_23, w_14_24, w_14_25, w_14_26, w_14_27, w_14_28, w_14_29, w_14_30, w_14_31, w_14_32, w_14_33, w_14_34, w_14_35, w_14_36, w_14_37, w_14_38, w_14_39, w_14_40, w_14_41, w_14_42, w_14_43, w_14_44, w_14_45;
    wire s_14_14, s_14_15, s_14_16, s_14_17, s_14_18, s_14_19, s_14_20, s_14_21, s_14_22, s_14_23, s_14_24, s_14_25, s_14_26, s_14_27, s_14_28, s_14_29, s_14_30, s_14_31, s_14_32, s_14_33, s_14_34, s_14_35, s_14_36, s_14_37, s_14_38, s_14_39, s_14_40, s_14_41, s_14_42, s_14_43, s_14_44, s_14_45;
    wire c_14_14, c_14_15, c_14_16, c_14_17, c_14_18, c_14_19, c_14_20, c_14_21, c_14_22, c_14_23, c_14_24, c_14_25, c_14_26, c_14_27, c_14_28, c_14_29, c_14_30, c_14_31, c_14_32, c_14_33, c_14_34, c_14_35, c_14_36, c_14_37, c_14_38, c_14_39, c_14_40, c_14_41, c_14_42, c_14_43, c_14_44, c_14_45;
    assign w_14_14 = data_operandA[0] & data_operandB[14];
    assign w_14_15 = data_operandA[1] & data_operandB[14];
    assign w_14_16 = data_operandA[2] & data_operandB[14];
    assign w_14_17 = data_operandA[3] & data_operandB[14];
    assign w_14_18 = data_operandA[4] & data_operandB[14];
    assign w_14_19 = data_operandA[5] & data_operandB[14];
    assign w_14_20 = data_operandA[6] & data_operandB[14];
    assign w_14_21 = data_operandA[7] & data_operandB[14];
    assign w_14_22 = data_operandA[8] & data_operandB[14];
    assign w_14_23 = data_operandA[9] & data_operandB[14];
    assign w_14_24 = data_operandA[10] & data_operandB[14];
    assign w_14_25 = data_operandA[11] & data_operandB[14];
    assign w_14_26 = data_operandA[12] & data_operandB[14];
    assign w_14_27 = data_operandA[13] & data_operandB[14];
    assign w_14_28 = data_operandA[14] & data_operandB[14];
    assign w_14_29 = data_operandA[15] & data_operandB[14];
    assign w_14_30 = data_operandA[16] & data_operandB[14];
    assign w_14_31 = data_operandA[17] & data_operandB[14];
    assign w_14_32 = data_operandA[18] & data_operandB[14];
    assign w_14_33 = data_operandA[19] & data_operandB[14];
    assign w_14_34 = data_operandA[20] & data_operandB[14];
    assign w_14_35 = data_operandA[21] & data_operandB[14];
    assign w_14_36 = data_operandA[22] & data_operandB[14];
    assign w_14_37 = data_operandA[23] & data_operandB[14];
    assign w_14_38 = data_operandA[24] & data_operandB[14];
    assign w_14_39 = data_operandA[25] & data_operandB[14];
    assign w_14_40 = data_operandA[26] & data_operandB[14];
    assign w_14_41 = data_operandA[27] & data_operandB[14];
    assign w_14_42 = data_operandA[28] & data_operandB[14];
    assign w_14_43 = data_operandA[29] & data_operandB[14];
    assign w_14_44 = data_operandA[30] & data_operandB[14];
    assign w_14_45 = ~(data_operandA[31] & data_operandB[14]);
    full_adder adder_14_14(.S(s_14_14), .Cout(c_14_14), .A(s_13_14), .B(w_14_14), .Cin(1'b0));
    full_adder adder_14_15(.S(s_14_15), .Cout(c_14_15), .A(s_13_15), .B(w_14_15), .Cin(c_14_14));
    full_adder adder_14_16(.S(s_14_16), .Cout(c_14_16), .A(s_13_16), .B(w_14_16), .Cin(c_14_15));
    full_adder adder_14_17(.S(s_14_17), .Cout(c_14_17), .A(s_13_17), .B(w_14_17), .Cin(c_14_16));
    full_adder adder_14_18(.S(s_14_18), .Cout(c_14_18), .A(s_13_18), .B(w_14_18), .Cin(c_14_17));
    full_adder adder_14_19(.S(s_14_19), .Cout(c_14_19), .A(s_13_19), .B(w_14_19), .Cin(c_14_18));
    full_adder adder_14_20(.S(s_14_20), .Cout(c_14_20), .A(s_13_20), .B(w_14_20), .Cin(c_14_19));
    full_adder adder_14_21(.S(s_14_21), .Cout(c_14_21), .A(s_13_21), .B(w_14_21), .Cin(c_14_20));
    full_adder adder_14_22(.S(s_14_22), .Cout(c_14_22), .A(s_13_22), .B(w_14_22), .Cin(c_14_21));
    full_adder adder_14_23(.S(s_14_23), .Cout(c_14_23), .A(s_13_23), .B(w_14_23), .Cin(c_14_22));
    full_adder adder_14_24(.S(s_14_24), .Cout(c_14_24), .A(s_13_24), .B(w_14_24), .Cin(c_14_23));
    full_adder adder_14_25(.S(s_14_25), .Cout(c_14_25), .A(s_13_25), .B(w_14_25), .Cin(c_14_24));
    full_adder adder_14_26(.S(s_14_26), .Cout(c_14_26), .A(s_13_26), .B(w_14_26), .Cin(c_14_25));
    full_adder adder_14_27(.S(s_14_27), .Cout(c_14_27), .A(s_13_27), .B(w_14_27), .Cin(c_14_26));
    full_adder adder_14_28(.S(s_14_28), .Cout(c_14_28), .A(s_13_28), .B(w_14_28), .Cin(c_14_27));
    full_adder adder_14_29(.S(s_14_29), .Cout(c_14_29), .A(s_13_29), .B(w_14_29), .Cin(c_14_28));
    full_adder adder_14_30(.S(s_14_30), .Cout(c_14_30), .A(s_13_30), .B(w_14_30), .Cin(c_14_29));
    full_adder adder_14_31(.S(s_14_31), .Cout(c_14_31), .A(s_13_31), .B(w_14_31), .Cin(c_14_30));
    full_adder adder_14_32(.S(s_14_32), .Cout(c_14_32), .A(s_13_32), .B(w_14_32), .Cin(c_14_31));
    full_adder adder_14_33(.S(s_14_33), .Cout(c_14_33), .A(s_13_33), .B(w_14_33), .Cin(c_14_32));
    full_adder adder_14_34(.S(s_14_34), .Cout(c_14_34), .A(s_13_34), .B(w_14_34), .Cin(c_14_33));
    full_adder adder_14_35(.S(s_14_35), .Cout(c_14_35), .A(s_13_35), .B(w_14_35), .Cin(c_14_34));
    full_adder adder_14_36(.S(s_14_36), .Cout(c_14_36), .A(s_13_36), .B(w_14_36), .Cin(c_14_35));
    full_adder adder_14_37(.S(s_14_37), .Cout(c_14_37), .A(s_13_37), .B(w_14_37), .Cin(c_14_36));
    full_adder adder_14_38(.S(s_14_38), .Cout(c_14_38), .A(s_13_38), .B(w_14_38), .Cin(c_14_37));
    full_adder adder_14_39(.S(s_14_39), .Cout(c_14_39), .A(s_13_39), .B(w_14_39), .Cin(c_14_38));
    full_adder adder_14_40(.S(s_14_40), .Cout(c_14_40), .A(s_13_40), .B(w_14_40), .Cin(c_14_39));
    full_adder adder_14_41(.S(s_14_41), .Cout(c_14_41), .A(s_13_41), .B(w_14_41), .Cin(c_14_40));
    full_adder adder_14_42(.S(s_14_42), .Cout(c_14_42), .A(s_13_42), .B(w_14_42), .Cin(c_14_41));
    full_adder adder_14_43(.S(s_14_43), .Cout(c_14_43), .A(s_13_43), .B(w_14_43), .Cin(c_14_42));
    full_adder adder_14_44(.S(s_14_44), .Cout(c_14_44), .A(s_13_44), .B(w_14_44), .Cin(c_14_43));
    full_adder adder_14_45(.S(s_14_45), .Cout(c_14_45), .A(c_13_44), .B(w_14_45), .Cin(c_14_44));
    assign result[14] = s_14_14;
    wire w_15_15, w_15_16, w_15_17, w_15_18, w_15_19, w_15_20, w_15_21, w_15_22, w_15_23, w_15_24, w_15_25, w_15_26, w_15_27, w_15_28, w_15_29, w_15_30, w_15_31, w_15_32, w_15_33, w_15_34, w_15_35, w_15_36, w_15_37, w_15_38, w_15_39, w_15_40, w_15_41, w_15_42, w_15_43, w_15_44, w_15_45, w_15_46;
    wire s_15_15, s_15_16, s_15_17, s_15_18, s_15_19, s_15_20, s_15_21, s_15_22, s_15_23, s_15_24, s_15_25, s_15_26, s_15_27, s_15_28, s_15_29, s_15_30, s_15_31, s_15_32, s_15_33, s_15_34, s_15_35, s_15_36, s_15_37, s_15_38, s_15_39, s_15_40, s_15_41, s_15_42, s_15_43, s_15_44, s_15_45, s_15_46;
    wire c_15_15, c_15_16, c_15_17, c_15_18, c_15_19, c_15_20, c_15_21, c_15_22, c_15_23, c_15_24, c_15_25, c_15_26, c_15_27, c_15_28, c_15_29, c_15_30, c_15_31, c_15_32, c_15_33, c_15_34, c_15_35, c_15_36, c_15_37, c_15_38, c_15_39, c_15_40, c_15_41, c_15_42, c_15_43, c_15_44, c_15_45, c_15_46;
    assign w_15_15 = data_operandA[0] & data_operandB[15];
    assign w_15_16 = data_operandA[1] & data_operandB[15];
    assign w_15_17 = data_operandA[2] & data_operandB[15];
    assign w_15_18 = data_operandA[3] & data_operandB[15];
    assign w_15_19 = data_operandA[4] & data_operandB[15];
    assign w_15_20 = data_operandA[5] & data_operandB[15];
    assign w_15_21 = data_operandA[6] & data_operandB[15];
    assign w_15_22 = data_operandA[7] & data_operandB[15];
    assign w_15_23 = data_operandA[8] & data_operandB[15];
    assign w_15_24 = data_operandA[9] & data_operandB[15];
    assign w_15_25 = data_operandA[10] & data_operandB[15];
    assign w_15_26 = data_operandA[11] & data_operandB[15];
    assign w_15_27 = data_operandA[12] & data_operandB[15];
    assign w_15_28 = data_operandA[13] & data_operandB[15];
    assign w_15_29 = data_operandA[14] & data_operandB[15];
    assign w_15_30 = data_operandA[15] & data_operandB[15];
    assign w_15_31 = data_operandA[16] & data_operandB[15];
    assign w_15_32 = data_operandA[17] & data_operandB[15];
    assign w_15_33 = data_operandA[18] & data_operandB[15];
    assign w_15_34 = data_operandA[19] & data_operandB[15];
    assign w_15_35 = data_operandA[20] & data_operandB[15];
    assign w_15_36 = data_operandA[21] & data_operandB[15];
    assign w_15_37 = data_operandA[22] & data_operandB[15];
    assign w_15_38 = data_operandA[23] & data_operandB[15];
    assign w_15_39 = data_operandA[24] & data_operandB[15];
    assign w_15_40 = data_operandA[25] & data_operandB[15];
    assign w_15_41 = data_operandA[26] & data_operandB[15];
    assign w_15_42 = data_operandA[27] & data_operandB[15];
    assign w_15_43 = data_operandA[28] & data_operandB[15];
    assign w_15_44 = data_operandA[29] & data_operandB[15];
    assign w_15_45 = data_operandA[30] & data_operandB[15];
    assign w_15_46 = ~(data_operandA[31] & data_operandB[15]);
    full_adder adder_15_15(.S(s_15_15), .Cout(c_15_15), .A(s_14_15), .B(w_15_15), .Cin(1'b0));
    full_adder adder_15_16(.S(s_15_16), .Cout(c_15_16), .A(s_14_16), .B(w_15_16), .Cin(c_15_15));
    full_adder adder_15_17(.S(s_15_17), .Cout(c_15_17), .A(s_14_17), .B(w_15_17), .Cin(c_15_16));
    full_adder adder_15_18(.S(s_15_18), .Cout(c_15_18), .A(s_14_18), .B(w_15_18), .Cin(c_15_17));
    full_adder adder_15_19(.S(s_15_19), .Cout(c_15_19), .A(s_14_19), .B(w_15_19), .Cin(c_15_18));
    full_adder adder_15_20(.S(s_15_20), .Cout(c_15_20), .A(s_14_20), .B(w_15_20), .Cin(c_15_19));
    full_adder adder_15_21(.S(s_15_21), .Cout(c_15_21), .A(s_14_21), .B(w_15_21), .Cin(c_15_20));
    full_adder adder_15_22(.S(s_15_22), .Cout(c_15_22), .A(s_14_22), .B(w_15_22), .Cin(c_15_21));
    full_adder adder_15_23(.S(s_15_23), .Cout(c_15_23), .A(s_14_23), .B(w_15_23), .Cin(c_15_22));
    full_adder adder_15_24(.S(s_15_24), .Cout(c_15_24), .A(s_14_24), .B(w_15_24), .Cin(c_15_23));
    full_adder adder_15_25(.S(s_15_25), .Cout(c_15_25), .A(s_14_25), .B(w_15_25), .Cin(c_15_24));
    full_adder adder_15_26(.S(s_15_26), .Cout(c_15_26), .A(s_14_26), .B(w_15_26), .Cin(c_15_25));
    full_adder adder_15_27(.S(s_15_27), .Cout(c_15_27), .A(s_14_27), .B(w_15_27), .Cin(c_15_26));
    full_adder adder_15_28(.S(s_15_28), .Cout(c_15_28), .A(s_14_28), .B(w_15_28), .Cin(c_15_27));
    full_adder adder_15_29(.S(s_15_29), .Cout(c_15_29), .A(s_14_29), .B(w_15_29), .Cin(c_15_28));
    full_adder adder_15_30(.S(s_15_30), .Cout(c_15_30), .A(s_14_30), .B(w_15_30), .Cin(c_15_29));
    full_adder adder_15_31(.S(s_15_31), .Cout(c_15_31), .A(s_14_31), .B(w_15_31), .Cin(c_15_30));
    full_adder adder_15_32(.S(s_15_32), .Cout(c_15_32), .A(s_14_32), .B(w_15_32), .Cin(c_15_31));
    full_adder adder_15_33(.S(s_15_33), .Cout(c_15_33), .A(s_14_33), .B(w_15_33), .Cin(c_15_32));
    full_adder adder_15_34(.S(s_15_34), .Cout(c_15_34), .A(s_14_34), .B(w_15_34), .Cin(c_15_33));
    full_adder adder_15_35(.S(s_15_35), .Cout(c_15_35), .A(s_14_35), .B(w_15_35), .Cin(c_15_34));
    full_adder adder_15_36(.S(s_15_36), .Cout(c_15_36), .A(s_14_36), .B(w_15_36), .Cin(c_15_35));
    full_adder adder_15_37(.S(s_15_37), .Cout(c_15_37), .A(s_14_37), .B(w_15_37), .Cin(c_15_36));
    full_adder adder_15_38(.S(s_15_38), .Cout(c_15_38), .A(s_14_38), .B(w_15_38), .Cin(c_15_37));
    full_adder adder_15_39(.S(s_15_39), .Cout(c_15_39), .A(s_14_39), .B(w_15_39), .Cin(c_15_38));
    full_adder adder_15_40(.S(s_15_40), .Cout(c_15_40), .A(s_14_40), .B(w_15_40), .Cin(c_15_39));
    full_adder adder_15_41(.S(s_15_41), .Cout(c_15_41), .A(s_14_41), .B(w_15_41), .Cin(c_15_40));
    full_adder adder_15_42(.S(s_15_42), .Cout(c_15_42), .A(s_14_42), .B(w_15_42), .Cin(c_15_41));
    full_adder adder_15_43(.S(s_15_43), .Cout(c_15_43), .A(s_14_43), .B(w_15_43), .Cin(c_15_42));
    full_adder adder_15_44(.S(s_15_44), .Cout(c_15_44), .A(s_14_44), .B(w_15_44), .Cin(c_15_43));
    full_adder adder_15_45(.S(s_15_45), .Cout(c_15_45), .A(s_14_45), .B(w_15_45), .Cin(c_15_44));
    full_adder adder_15_46(.S(s_15_46), .Cout(c_15_46), .A(c_14_45), .B(w_15_46), .Cin(c_15_45));
    assign result[15] = s_15_15;
    wire w_16_16, w_16_17, w_16_18, w_16_19, w_16_20, w_16_21, w_16_22, w_16_23, w_16_24, w_16_25, w_16_26, w_16_27, w_16_28, w_16_29, w_16_30, w_16_31, w_16_32, w_16_33, w_16_34, w_16_35, w_16_36, w_16_37, w_16_38, w_16_39, w_16_40, w_16_41, w_16_42, w_16_43, w_16_44, w_16_45, w_16_46, w_16_47;
    wire s_16_16, s_16_17, s_16_18, s_16_19, s_16_20, s_16_21, s_16_22, s_16_23, s_16_24, s_16_25, s_16_26, s_16_27, s_16_28, s_16_29, s_16_30, s_16_31, s_16_32, s_16_33, s_16_34, s_16_35, s_16_36, s_16_37, s_16_38, s_16_39, s_16_40, s_16_41, s_16_42, s_16_43, s_16_44, s_16_45, s_16_46, s_16_47;
    wire c_16_16, c_16_17, c_16_18, c_16_19, c_16_20, c_16_21, c_16_22, c_16_23, c_16_24, c_16_25, c_16_26, c_16_27, c_16_28, c_16_29, c_16_30, c_16_31, c_16_32, c_16_33, c_16_34, c_16_35, c_16_36, c_16_37, c_16_38, c_16_39, c_16_40, c_16_41, c_16_42, c_16_43, c_16_44, c_16_45, c_16_46, c_16_47;
    assign w_16_16 = data_operandA[0] & data_operandB[16];
    assign w_16_17 = data_operandA[1] & data_operandB[16];
    assign w_16_18 = data_operandA[2] & data_operandB[16];
    assign w_16_19 = data_operandA[3] & data_operandB[16];
    assign w_16_20 = data_operandA[4] & data_operandB[16];
    assign w_16_21 = data_operandA[5] & data_operandB[16];
    assign w_16_22 = data_operandA[6] & data_operandB[16];
    assign w_16_23 = data_operandA[7] & data_operandB[16];
    assign w_16_24 = data_operandA[8] & data_operandB[16];
    assign w_16_25 = data_operandA[9] & data_operandB[16];
    assign w_16_26 = data_operandA[10] & data_operandB[16];
    assign w_16_27 = data_operandA[11] & data_operandB[16];
    assign w_16_28 = data_operandA[12] & data_operandB[16];
    assign w_16_29 = data_operandA[13] & data_operandB[16];
    assign w_16_30 = data_operandA[14] & data_operandB[16];
    assign w_16_31 = data_operandA[15] & data_operandB[16];
    assign w_16_32 = data_operandA[16] & data_operandB[16];
    assign w_16_33 = data_operandA[17] & data_operandB[16];
    assign w_16_34 = data_operandA[18] & data_operandB[16];
    assign w_16_35 = data_operandA[19] & data_operandB[16];
    assign w_16_36 = data_operandA[20] & data_operandB[16];
    assign w_16_37 = data_operandA[21] & data_operandB[16];
    assign w_16_38 = data_operandA[22] & data_operandB[16];
    assign w_16_39 = data_operandA[23] & data_operandB[16];
    assign w_16_40 = data_operandA[24] & data_operandB[16];
    assign w_16_41 = data_operandA[25] & data_operandB[16];
    assign w_16_42 = data_operandA[26] & data_operandB[16];
    assign w_16_43 = data_operandA[27] & data_operandB[16];
    assign w_16_44 = data_operandA[28] & data_operandB[16];
    assign w_16_45 = data_operandA[29] & data_operandB[16];
    assign w_16_46 = data_operandA[30] & data_operandB[16];
    assign w_16_47 = ~(data_operandA[31] & data_operandB[16]);
    full_adder adder_16_16(.S(s_16_16), .Cout(c_16_16), .A(s_15_16), .B(w_16_16), .Cin(1'b0));
    full_adder adder_16_17(.S(s_16_17), .Cout(c_16_17), .A(s_15_17), .B(w_16_17), .Cin(c_16_16));
    full_adder adder_16_18(.S(s_16_18), .Cout(c_16_18), .A(s_15_18), .B(w_16_18), .Cin(c_16_17));
    full_adder adder_16_19(.S(s_16_19), .Cout(c_16_19), .A(s_15_19), .B(w_16_19), .Cin(c_16_18));
    full_adder adder_16_20(.S(s_16_20), .Cout(c_16_20), .A(s_15_20), .B(w_16_20), .Cin(c_16_19));
    full_adder adder_16_21(.S(s_16_21), .Cout(c_16_21), .A(s_15_21), .B(w_16_21), .Cin(c_16_20));
    full_adder adder_16_22(.S(s_16_22), .Cout(c_16_22), .A(s_15_22), .B(w_16_22), .Cin(c_16_21));
    full_adder adder_16_23(.S(s_16_23), .Cout(c_16_23), .A(s_15_23), .B(w_16_23), .Cin(c_16_22));
    full_adder adder_16_24(.S(s_16_24), .Cout(c_16_24), .A(s_15_24), .B(w_16_24), .Cin(c_16_23));
    full_adder adder_16_25(.S(s_16_25), .Cout(c_16_25), .A(s_15_25), .B(w_16_25), .Cin(c_16_24));
    full_adder adder_16_26(.S(s_16_26), .Cout(c_16_26), .A(s_15_26), .B(w_16_26), .Cin(c_16_25));
    full_adder adder_16_27(.S(s_16_27), .Cout(c_16_27), .A(s_15_27), .B(w_16_27), .Cin(c_16_26));
    full_adder adder_16_28(.S(s_16_28), .Cout(c_16_28), .A(s_15_28), .B(w_16_28), .Cin(c_16_27));
    full_adder adder_16_29(.S(s_16_29), .Cout(c_16_29), .A(s_15_29), .B(w_16_29), .Cin(c_16_28));
    full_adder adder_16_30(.S(s_16_30), .Cout(c_16_30), .A(s_15_30), .B(w_16_30), .Cin(c_16_29));
    full_adder adder_16_31(.S(s_16_31), .Cout(c_16_31), .A(s_15_31), .B(w_16_31), .Cin(c_16_30));
    full_adder adder_16_32(.S(s_16_32), .Cout(c_16_32), .A(s_15_32), .B(w_16_32), .Cin(c_16_31));
    full_adder adder_16_33(.S(s_16_33), .Cout(c_16_33), .A(s_15_33), .B(w_16_33), .Cin(c_16_32));
    full_adder adder_16_34(.S(s_16_34), .Cout(c_16_34), .A(s_15_34), .B(w_16_34), .Cin(c_16_33));
    full_adder adder_16_35(.S(s_16_35), .Cout(c_16_35), .A(s_15_35), .B(w_16_35), .Cin(c_16_34));
    full_adder adder_16_36(.S(s_16_36), .Cout(c_16_36), .A(s_15_36), .B(w_16_36), .Cin(c_16_35));
    full_adder adder_16_37(.S(s_16_37), .Cout(c_16_37), .A(s_15_37), .B(w_16_37), .Cin(c_16_36));
    full_adder adder_16_38(.S(s_16_38), .Cout(c_16_38), .A(s_15_38), .B(w_16_38), .Cin(c_16_37));
    full_adder adder_16_39(.S(s_16_39), .Cout(c_16_39), .A(s_15_39), .B(w_16_39), .Cin(c_16_38));
    full_adder adder_16_40(.S(s_16_40), .Cout(c_16_40), .A(s_15_40), .B(w_16_40), .Cin(c_16_39));
    full_adder adder_16_41(.S(s_16_41), .Cout(c_16_41), .A(s_15_41), .B(w_16_41), .Cin(c_16_40));
    full_adder adder_16_42(.S(s_16_42), .Cout(c_16_42), .A(s_15_42), .B(w_16_42), .Cin(c_16_41));
    full_adder adder_16_43(.S(s_16_43), .Cout(c_16_43), .A(s_15_43), .B(w_16_43), .Cin(c_16_42));
    full_adder adder_16_44(.S(s_16_44), .Cout(c_16_44), .A(s_15_44), .B(w_16_44), .Cin(c_16_43));
    full_adder adder_16_45(.S(s_16_45), .Cout(c_16_45), .A(s_15_45), .B(w_16_45), .Cin(c_16_44));
    full_adder adder_16_46(.S(s_16_46), .Cout(c_16_46), .A(s_15_46), .B(w_16_46), .Cin(c_16_45));
    full_adder adder_16_47(.S(s_16_47), .Cout(c_16_47), .A(c_15_46), .B(w_16_47), .Cin(c_16_46));
    assign result[16] = s_16_16;
    wire w_17_17, w_17_18, w_17_19, w_17_20, w_17_21, w_17_22, w_17_23, w_17_24, w_17_25, w_17_26, w_17_27, w_17_28, w_17_29, w_17_30, w_17_31, w_17_32, w_17_33, w_17_34, w_17_35, w_17_36, w_17_37, w_17_38, w_17_39, w_17_40, w_17_41, w_17_42, w_17_43, w_17_44, w_17_45, w_17_46, w_17_47, w_17_48;
    wire s_17_17, s_17_18, s_17_19, s_17_20, s_17_21, s_17_22, s_17_23, s_17_24, s_17_25, s_17_26, s_17_27, s_17_28, s_17_29, s_17_30, s_17_31, s_17_32, s_17_33, s_17_34, s_17_35, s_17_36, s_17_37, s_17_38, s_17_39, s_17_40, s_17_41, s_17_42, s_17_43, s_17_44, s_17_45, s_17_46, s_17_47, s_17_48;
    wire c_17_17, c_17_18, c_17_19, c_17_20, c_17_21, c_17_22, c_17_23, c_17_24, c_17_25, c_17_26, c_17_27, c_17_28, c_17_29, c_17_30, c_17_31, c_17_32, c_17_33, c_17_34, c_17_35, c_17_36, c_17_37, c_17_38, c_17_39, c_17_40, c_17_41, c_17_42, c_17_43, c_17_44, c_17_45, c_17_46, c_17_47, c_17_48;
    assign w_17_17 = data_operandA[0] & data_operandB[17];
    assign w_17_18 = data_operandA[1] & data_operandB[17];
    assign w_17_19 = data_operandA[2] & data_operandB[17];
    assign w_17_20 = data_operandA[3] & data_operandB[17];
    assign w_17_21 = data_operandA[4] & data_operandB[17];
    assign w_17_22 = data_operandA[5] & data_operandB[17];
    assign w_17_23 = data_operandA[6] & data_operandB[17];
    assign w_17_24 = data_operandA[7] & data_operandB[17];
    assign w_17_25 = data_operandA[8] & data_operandB[17];
    assign w_17_26 = data_operandA[9] & data_operandB[17];
    assign w_17_27 = data_operandA[10] & data_operandB[17];
    assign w_17_28 = data_operandA[11] & data_operandB[17];
    assign w_17_29 = data_operandA[12] & data_operandB[17];
    assign w_17_30 = data_operandA[13] & data_operandB[17];
    assign w_17_31 = data_operandA[14] & data_operandB[17];
    assign w_17_32 = data_operandA[15] & data_operandB[17];
    assign w_17_33 = data_operandA[16] & data_operandB[17];
    assign w_17_34 = data_operandA[17] & data_operandB[17];
    assign w_17_35 = data_operandA[18] & data_operandB[17];
    assign w_17_36 = data_operandA[19] & data_operandB[17];
    assign w_17_37 = data_operandA[20] & data_operandB[17];
    assign w_17_38 = data_operandA[21] & data_operandB[17];
    assign w_17_39 = data_operandA[22] & data_operandB[17];
    assign w_17_40 = data_operandA[23] & data_operandB[17];
    assign w_17_41 = data_operandA[24] & data_operandB[17];
    assign w_17_42 = data_operandA[25] & data_operandB[17];
    assign w_17_43 = data_operandA[26] & data_operandB[17];
    assign w_17_44 = data_operandA[27] & data_operandB[17];
    assign w_17_45 = data_operandA[28] & data_operandB[17];
    assign w_17_46 = data_operandA[29] & data_operandB[17];
    assign w_17_47 = data_operandA[30] & data_operandB[17];
    assign w_17_48 = ~(data_operandA[31] & data_operandB[17]);
    full_adder adder_17_17(.S(s_17_17), .Cout(c_17_17), .A(s_16_17), .B(w_17_17), .Cin(1'b0));
    full_adder adder_17_18(.S(s_17_18), .Cout(c_17_18), .A(s_16_18), .B(w_17_18), .Cin(c_17_17));
    full_adder adder_17_19(.S(s_17_19), .Cout(c_17_19), .A(s_16_19), .B(w_17_19), .Cin(c_17_18));
    full_adder adder_17_20(.S(s_17_20), .Cout(c_17_20), .A(s_16_20), .B(w_17_20), .Cin(c_17_19));
    full_adder adder_17_21(.S(s_17_21), .Cout(c_17_21), .A(s_16_21), .B(w_17_21), .Cin(c_17_20));
    full_adder adder_17_22(.S(s_17_22), .Cout(c_17_22), .A(s_16_22), .B(w_17_22), .Cin(c_17_21));
    full_adder adder_17_23(.S(s_17_23), .Cout(c_17_23), .A(s_16_23), .B(w_17_23), .Cin(c_17_22));
    full_adder adder_17_24(.S(s_17_24), .Cout(c_17_24), .A(s_16_24), .B(w_17_24), .Cin(c_17_23));
    full_adder adder_17_25(.S(s_17_25), .Cout(c_17_25), .A(s_16_25), .B(w_17_25), .Cin(c_17_24));
    full_adder adder_17_26(.S(s_17_26), .Cout(c_17_26), .A(s_16_26), .B(w_17_26), .Cin(c_17_25));
    full_adder adder_17_27(.S(s_17_27), .Cout(c_17_27), .A(s_16_27), .B(w_17_27), .Cin(c_17_26));
    full_adder adder_17_28(.S(s_17_28), .Cout(c_17_28), .A(s_16_28), .B(w_17_28), .Cin(c_17_27));
    full_adder adder_17_29(.S(s_17_29), .Cout(c_17_29), .A(s_16_29), .B(w_17_29), .Cin(c_17_28));
    full_adder adder_17_30(.S(s_17_30), .Cout(c_17_30), .A(s_16_30), .B(w_17_30), .Cin(c_17_29));
    full_adder adder_17_31(.S(s_17_31), .Cout(c_17_31), .A(s_16_31), .B(w_17_31), .Cin(c_17_30));
    full_adder adder_17_32(.S(s_17_32), .Cout(c_17_32), .A(s_16_32), .B(w_17_32), .Cin(c_17_31));
    full_adder adder_17_33(.S(s_17_33), .Cout(c_17_33), .A(s_16_33), .B(w_17_33), .Cin(c_17_32));
    full_adder adder_17_34(.S(s_17_34), .Cout(c_17_34), .A(s_16_34), .B(w_17_34), .Cin(c_17_33));
    full_adder adder_17_35(.S(s_17_35), .Cout(c_17_35), .A(s_16_35), .B(w_17_35), .Cin(c_17_34));
    full_adder adder_17_36(.S(s_17_36), .Cout(c_17_36), .A(s_16_36), .B(w_17_36), .Cin(c_17_35));
    full_adder adder_17_37(.S(s_17_37), .Cout(c_17_37), .A(s_16_37), .B(w_17_37), .Cin(c_17_36));
    full_adder adder_17_38(.S(s_17_38), .Cout(c_17_38), .A(s_16_38), .B(w_17_38), .Cin(c_17_37));
    full_adder adder_17_39(.S(s_17_39), .Cout(c_17_39), .A(s_16_39), .B(w_17_39), .Cin(c_17_38));
    full_adder adder_17_40(.S(s_17_40), .Cout(c_17_40), .A(s_16_40), .B(w_17_40), .Cin(c_17_39));
    full_adder adder_17_41(.S(s_17_41), .Cout(c_17_41), .A(s_16_41), .B(w_17_41), .Cin(c_17_40));
    full_adder adder_17_42(.S(s_17_42), .Cout(c_17_42), .A(s_16_42), .B(w_17_42), .Cin(c_17_41));
    full_adder adder_17_43(.S(s_17_43), .Cout(c_17_43), .A(s_16_43), .B(w_17_43), .Cin(c_17_42));
    full_adder adder_17_44(.S(s_17_44), .Cout(c_17_44), .A(s_16_44), .B(w_17_44), .Cin(c_17_43));
    full_adder adder_17_45(.S(s_17_45), .Cout(c_17_45), .A(s_16_45), .B(w_17_45), .Cin(c_17_44));
    full_adder adder_17_46(.S(s_17_46), .Cout(c_17_46), .A(s_16_46), .B(w_17_46), .Cin(c_17_45));
    full_adder adder_17_47(.S(s_17_47), .Cout(c_17_47), .A(s_16_47), .B(w_17_47), .Cin(c_17_46));
    full_adder adder_17_48(.S(s_17_48), .Cout(c_17_48), .A(c_16_47), .B(w_17_48), .Cin(c_17_47));
    assign result[17] = s_17_17;
    wire w_18_18, w_18_19, w_18_20, w_18_21, w_18_22, w_18_23, w_18_24, w_18_25, w_18_26, w_18_27, w_18_28, w_18_29, w_18_30, w_18_31, w_18_32, w_18_33, w_18_34, w_18_35, w_18_36, w_18_37, w_18_38, w_18_39, w_18_40, w_18_41, w_18_42, w_18_43, w_18_44, w_18_45, w_18_46, w_18_47, w_18_48, w_18_49;
    wire s_18_18, s_18_19, s_18_20, s_18_21, s_18_22, s_18_23, s_18_24, s_18_25, s_18_26, s_18_27, s_18_28, s_18_29, s_18_30, s_18_31, s_18_32, s_18_33, s_18_34, s_18_35, s_18_36, s_18_37, s_18_38, s_18_39, s_18_40, s_18_41, s_18_42, s_18_43, s_18_44, s_18_45, s_18_46, s_18_47, s_18_48, s_18_49;
    wire c_18_18, c_18_19, c_18_20, c_18_21, c_18_22, c_18_23, c_18_24, c_18_25, c_18_26, c_18_27, c_18_28, c_18_29, c_18_30, c_18_31, c_18_32, c_18_33, c_18_34, c_18_35, c_18_36, c_18_37, c_18_38, c_18_39, c_18_40, c_18_41, c_18_42, c_18_43, c_18_44, c_18_45, c_18_46, c_18_47, c_18_48, c_18_49;
    assign w_18_18 = data_operandA[0] & data_operandB[18];
    assign w_18_19 = data_operandA[1] & data_operandB[18];
    assign w_18_20 = data_operandA[2] & data_operandB[18];
    assign w_18_21 = data_operandA[3] & data_operandB[18];
    assign w_18_22 = data_operandA[4] & data_operandB[18];
    assign w_18_23 = data_operandA[5] & data_operandB[18];
    assign w_18_24 = data_operandA[6] & data_operandB[18];
    assign w_18_25 = data_operandA[7] & data_operandB[18];
    assign w_18_26 = data_operandA[8] & data_operandB[18];
    assign w_18_27 = data_operandA[9] & data_operandB[18];
    assign w_18_28 = data_operandA[10] & data_operandB[18];
    assign w_18_29 = data_operandA[11] & data_operandB[18];
    assign w_18_30 = data_operandA[12] & data_operandB[18];
    assign w_18_31 = data_operandA[13] & data_operandB[18];
    assign w_18_32 = data_operandA[14] & data_operandB[18];
    assign w_18_33 = data_operandA[15] & data_operandB[18];
    assign w_18_34 = data_operandA[16] & data_operandB[18];
    assign w_18_35 = data_operandA[17] & data_operandB[18];
    assign w_18_36 = data_operandA[18] & data_operandB[18];
    assign w_18_37 = data_operandA[19] & data_operandB[18];
    assign w_18_38 = data_operandA[20] & data_operandB[18];
    assign w_18_39 = data_operandA[21] & data_operandB[18];
    assign w_18_40 = data_operandA[22] & data_operandB[18];
    assign w_18_41 = data_operandA[23] & data_operandB[18];
    assign w_18_42 = data_operandA[24] & data_operandB[18];
    assign w_18_43 = data_operandA[25] & data_operandB[18];
    assign w_18_44 = data_operandA[26] & data_operandB[18];
    assign w_18_45 = data_operandA[27] & data_operandB[18];
    assign w_18_46 = data_operandA[28] & data_operandB[18];
    assign w_18_47 = data_operandA[29] & data_operandB[18];
    assign w_18_48 = data_operandA[30] & data_operandB[18];
    assign w_18_49 = ~(data_operandA[31] & data_operandB[18]);
    full_adder adder_18_18(.S(s_18_18), .Cout(c_18_18), .A(s_17_18), .B(w_18_18), .Cin(1'b0));
    full_adder adder_18_19(.S(s_18_19), .Cout(c_18_19), .A(s_17_19), .B(w_18_19), .Cin(c_18_18));
    full_adder adder_18_20(.S(s_18_20), .Cout(c_18_20), .A(s_17_20), .B(w_18_20), .Cin(c_18_19));
    full_adder adder_18_21(.S(s_18_21), .Cout(c_18_21), .A(s_17_21), .B(w_18_21), .Cin(c_18_20));
    full_adder adder_18_22(.S(s_18_22), .Cout(c_18_22), .A(s_17_22), .B(w_18_22), .Cin(c_18_21));
    full_adder adder_18_23(.S(s_18_23), .Cout(c_18_23), .A(s_17_23), .B(w_18_23), .Cin(c_18_22));
    full_adder adder_18_24(.S(s_18_24), .Cout(c_18_24), .A(s_17_24), .B(w_18_24), .Cin(c_18_23));
    full_adder adder_18_25(.S(s_18_25), .Cout(c_18_25), .A(s_17_25), .B(w_18_25), .Cin(c_18_24));
    full_adder adder_18_26(.S(s_18_26), .Cout(c_18_26), .A(s_17_26), .B(w_18_26), .Cin(c_18_25));
    full_adder adder_18_27(.S(s_18_27), .Cout(c_18_27), .A(s_17_27), .B(w_18_27), .Cin(c_18_26));
    full_adder adder_18_28(.S(s_18_28), .Cout(c_18_28), .A(s_17_28), .B(w_18_28), .Cin(c_18_27));
    full_adder adder_18_29(.S(s_18_29), .Cout(c_18_29), .A(s_17_29), .B(w_18_29), .Cin(c_18_28));
    full_adder adder_18_30(.S(s_18_30), .Cout(c_18_30), .A(s_17_30), .B(w_18_30), .Cin(c_18_29));
    full_adder adder_18_31(.S(s_18_31), .Cout(c_18_31), .A(s_17_31), .B(w_18_31), .Cin(c_18_30));
    full_adder adder_18_32(.S(s_18_32), .Cout(c_18_32), .A(s_17_32), .B(w_18_32), .Cin(c_18_31));
    full_adder adder_18_33(.S(s_18_33), .Cout(c_18_33), .A(s_17_33), .B(w_18_33), .Cin(c_18_32));
    full_adder adder_18_34(.S(s_18_34), .Cout(c_18_34), .A(s_17_34), .B(w_18_34), .Cin(c_18_33));
    full_adder adder_18_35(.S(s_18_35), .Cout(c_18_35), .A(s_17_35), .B(w_18_35), .Cin(c_18_34));
    full_adder adder_18_36(.S(s_18_36), .Cout(c_18_36), .A(s_17_36), .B(w_18_36), .Cin(c_18_35));
    full_adder adder_18_37(.S(s_18_37), .Cout(c_18_37), .A(s_17_37), .B(w_18_37), .Cin(c_18_36));
    full_adder adder_18_38(.S(s_18_38), .Cout(c_18_38), .A(s_17_38), .B(w_18_38), .Cin(c_18_37));
    full_adder adder_18_39(.S(s_18_39), .Cout(c_18_39), .A(s_17_39), .B(w_18_39), .Cin(c_18_38));
    full_adder adder_18_40(.S(s_18_40), .Cout(c_18_40), .A(s_17_40), .B(w_18_40), .Cin(c_18_39));
    full_adder adder_18_41(.S(s_18_41), .Cout(c_18_41), .A(s_17_41), .B(w_18_41), .Cin(c_18_40));
    full_adder adder_18_42(.S(s_18_42), .Cout(c_18_42), .A(s_17_42), .B(w_18_42), .Cin(c_18_41));
    full_adder adder_18_43(.S(s_18_43), .Cout(c_18_43), .A(s_17_43), .B(w_18_43), .Cin(c_18_42));
    full_adder adder_18_44(.S(s_18_44), .Cout(c_18_44), .A(s_17_44), .B(w_18_44), .Cin(c_18_43));
    full_adder adder_18_45(.S(s_18_45), .Cout(c_18_45), .A(s_17_45), .B(w_18_45), .Cin(c_18_44));
    full_adder adder_18_46(.S(s_18_46), .Cout(c_18_46), .A(s_17_46), .B(w_18_46), .Cin(c_18_45));
    full_adder adder_18_47(.S(s_18_47), .Cout(c_18_47), .A(s_17_47), .B(w_18_47), .Cin(c_18_46));
    full_adder adder_18_48(.S(s_18_48), .Cout(c_18_48), .A(s_17_48), .B(w_18_48), .Cin(c_18_47));
    full_adder adder_18_49(.S(s_18_49), .Cout(c_18_49), .A(c_17_48), .B(w_18_49), .Cin(c_18_48));
    assign result[18] = s_18_18;
    wire w_19_19, w_19_20, w_19_21, w_19_22, w_19_23, w_19_24, w_19_25, w_19_26, w_19_27, w_19_28, w_19_29, w_19_30, w_19_31, w_19_32, w_19_33, w_19_34, w_19_35, w_19_36, w_19_37, w_19_38, w_19_39, w_19_40, w_19_41, w_19_42, w_19_43, w_19_44, w_19_45, w_19_46, w_19_47, w_19_48, w_19_49, w_19_50;
    wire s_19_19, s_19_20, s_19_21, s_19_22, s_19_23, s_19_24, s_19_25, s_19_26, s_19_27, s_19_28, s_19_29, s_19_30, s_19_31, s_19_32, s_19_33, s_19_34, s_19_35, s_19_36, s_19_37, s_19_38, s_19_39, s_19_40, s_19_41, s_19_42, s_19_43, s_19_44, s_19_45, s_19_46, s_19_47, s_19_48, s_19_49, s_19_50;
    wire c_19_19, c_19_20, c_19_21, c_19_22, c_19_23, c_19_24, c_19_25, c_19_26, c_19_27, c_19_28, c_19_29, c_19_30, c_19_31, c_19_32, c_19_33, c_19_34, c_19_35, c_19_36, c_19_37, c_19_38, c_19_39, c_19_40, c_19_41, c_19_42, c_19_43, c_19_44, c_19_45, c_19_46, c_19_47, c_19_48, c_19_49, c_19_50;
    assign w_19_19 = data_operandA[0] & data_operandB[19];
    assign w_19_20 = data_operandA[1] & data_operandB[19];
    assign w_19_21 = data_operandA[2] & data_operandB[19];
    assign w_19_22 = data_operandA[3] & data_operandB[19];
    assign w_19_23 = data_operandA[4] & data_operandB[19];
    assign w_19_24 = data_operandA[5] & data_operandB[19];
    assign w_19_25 = data_operandA[6] & data_operandB[19];
    assign w_19_26 = data_operandA[7] & data_operandB[19];
    assign w_19_27 = data_operandA[8] & data_operandB[19];
    assign w_19_28 = data_operandA[9] & data_operandB[19];
    assign w_19_29 = data_operandA[10] & data_operandB[19];
    assign w_19_30 = data_operandA[11] & data_operandB[19];
    assign w_19_31 = data_operandA[12] & data_operandB[19];
    assign w_19_32 = data_operandA[13] & data_operandB[19];
    assign w_19_33 = data_operandA[14] & data_operandB[19];
    assign w_19_34 = data_operandA[15] & data_operandB[19];
    assign w_19_35 = data_operandA[16] & data_operandB[19];
    assign w_19_36 = data_operandA[17] & data_operandB[19];
    assign w_19_37 = data_operandA[18] & data_operandB[19];
    assign w_19_38 = data_operandA[19] & data_operandB[19];
    assign w_19_39 = data_operandA[20] & data_operandB[19];
    assign w_19_40 = data_operandA[21] & data_operandB[19];
    assign w_19_41 = data_operandA[22] & data_operandB[19];
    assign w_19_42 = data_operandA[23] & data_operandB[19];
    assign w_19_43 = data_operandA[24] & data_operandB[19];
    assign w_19_44 = data_operandA[25] & data_operandB[19];
    assign w_19_45 = data_operandA[26] & data_operandB[19];
    assign w_19_46 = data_operandA[27] & data_operandB[19];
    assign w_19_47 = data_operandA[28] & data_operandB[19];
    assign w_19_48 = data_operandA[29] & data_operandB[19];
    assign w_19_49 = data_operandA[30] & data_operandB[19];
    assign w_19_50 = ~(data_operandA[31] & data_operandB[19]);
    full_adder adder_19_19(.S(s_19_19), .Cout(c_19_19), .A(s_18_19), .B(w_19_19), .Cin(1'b0));
    full_adder adder_19_20(.S(s_19_20), .Cout(c_19_20), .A(s_18_20), .B(w_19_20), .Cin(c_19_19));
    full_adder adder_19_21(.S(s_19_21), .Cout(c_19_21), .A(s_18_21), .B(w_19_21), .Cin(c_19_20));
    full_adder adder_19_22(.S(s_19_22), .Cout(c_19_22), .A(s_18_22), .B(w_19_22), .Cin(c_19_21));
    full_adder adder_19_23(.S(s_19_23), .Cout(c_19_23), .A(s_18_23), .B(w_19_23), .Cin(c_19_22));
    full_adder adder_19_24(.S(s_19_24), .Cout(c_19_24), .A(s_18_24), .B(w_19_24), .Cin(c_19_23));
    full_adder adder_19_25(.S(s_19_25), .Cout(c_19_25), .A(s_18_25), .B(w_19_25), .Cin(c_19_24));
    full_adder adder_19_26(.S(s_19_26), .Cout(c_19_26), .A(s_18_26), .B(w_19_26), .Cin(c_19_25));
    full_adder adder_19_27(.S(s_19_27), .Cout(c_19_27), .A(s_18_27), .B(w_19_27), .Cin(c_19_26));
    full_adder adder_19_28(.S(s_19_28), .Cout(c_19_28), .A(s_18_28), .B(w_19_28), .Cin(c_19_27));
    full_adder adder_19_29(.S(s_19_29), .Cout(c_19_29), .A(s_18_29), .B(w_19_29), .Cin(c_19_28));
    full_adder adder_19_30(.S(s_19_30), .Cout(c_19_30), .A(s_18_30), .B(w_19_30), .Cin(c_19_29));
    full_adder adder_19_31(.S(s_19_31), .Cout(c_19_31), .A(s_18_31), .B(w_19_31), .Cin(c_19_30));
    full_adder adder_19_32(.S(s_19_32), .Cout(c_19_32), .A(s_18_32), .B(w_19_32), .Cin(c_19_31));
    full_adder adder_19_33(.S(s_19_33), .Cout(c_19_33), .A(s_18_33), .B(w_19_33), .Cin(c_19_32));
    full_adder adder_19_34(.S(s_19_34), .Cout(c_19_34), .A(s_18_34), .B(w_19_34), .Cin(c_19_33));
    full_adder adder_19_35(.S(s_19_35), .Cout(c_19_35), .A(s_18_35), .B(w_19_35), .Cin(c_19_34));
    full_adder adder_19_36(.S(s_19_36), .Cout(c_19_36), .A(s_18_36), .B(w_19_36), .Cin(c_19_35));
    full_adder adder_19_37(.S(s_19_37), .Cout(c_19_37), .A(s_18_37), .B(w_19_37), .Cin(c_19_36));
    full_adder adder_19_38(.S(s_19_38), .Cout(c_19_38), .A(s_18_38), .B(w_19_38), .Cin(c_19_37));
    full_adder adder_19_39(.S(s_19_39), .Cout(c_19_39), .A(s_18_39), .B(w_19_39), .Cin(c_19_38));
    full_adder adder_19_40(.S(s_19_40), .Cout(c_19_40), .A(s_18_40), .B(w_19_40), .Cin(c_19_39));
    full_adder adder_19_41(.S(s_19_41), .Cout(c_19_41), .A(s_18_41), .B(w_19_41), .Cin(c_19_40));
    full_adder adder_19_42(.S(s_19_42), .Cout(c_19_42), .A(s_18_42), .B(w_19_42), .Cin(c_19_41));
    full_adder adder_19_43(.S(s_19_43), .Cout(c_19_43), .A(s_18_43), .B(w_19_43), .Cin(c_19_42));
    full_adder adder_19_44(.S(s_19_44), .Cout(c_19_44), .A(s_18_44), .B(w_19_44), .Cin(c_19_43));
    full_adder adder_19_45(.S(s_19_45), .Cout(c_19_45), .A(s_18_45), .B(w_19_45), .Cin(c_19_44));
    full_adder adder_19_46(.S(s_19_46), .Cout(c_19_46), .A(s_18_46), .B(w_19_46), .Cin(c_19_45));
    full_adder adder_19_47(.S(s_19_47), .Cout(c_19_47), .A(s_18_47), .B(w_19_47), .Cin(c_19_46));
    full_adder adder_19_48(.S(s_19_48), .Cout(c_19_48), .A(s_18_48), .B(w_19_48), .Cin(c_19_47));
    full_adder adder_19_49(.S(s_19_49), .Cout(c_19_49), .A(s_18_49), .B(w_19_49), .Cin(c_19_48));
    full_adder adder_19_50(.S(s_19_50), .Cout(c_19_50), .A(c_18_49), .B(w_19_50), .Cin(c_19_49));
    assign result[19] = s_19_19;
    wire w_20_20, w_20_21, w_20_22, w_20_23, w_20_24, w_20_25, w_20_26, w_20_27, w_20_28, w_20_29, w_20_30, w_20_31, w_20_32, w_20_33, w_20_34, w_20_35, w_20_36, w_20_37, w_20_38, w_20_39, w_20_40, w_20_41, w_20_42, w_20_43, w_20_44, w_20_45, w_20_46, w_20_47, w_20_48, w_20_49, w_20_50, w_20_51;
    wire s_20_20, s_20_21, s_20_22, s_20_23, s_20_24, s_20_25, s_20_26, s_20_27, s_20_28, s_20_29, s_20_30, s_20_31, s_20_32, s_20_33, s_20_34, s_20_35, s_20_36, s_20_37, s_20_38, s_20_39, s_20_40, s_20_41, s_20_42, s_20_43, s_20_44, s_20_45, s_20_46, s_20_47, s_20_48, s_20_49, s_20_50, s_20_51;
    wire c_20_20, c_20_21, c_20_22, c_20_23, c_20_24, c_20_25, c_20_26, c_20_27, c_20_28, c_20_29, c_20_30, c_20_31, c_20_32, c_20_33, c_20_34, c_20_35, c_20_36, c_20_37, c_20_38, c_20_39, c_20_40, c_20_41, c_20_42, c_20_43, c_20_44, c_20_45, c_20_46, c_20_47, c_20_48, c_20_49, c_20_50, c_20_51;
    assign w_20_20 = data_operandA[0] & data_operandB[20];
    assign w_20_21 = data_operandA[1] & data_operandB[20];
    assign w_20_22 = data_operandA[2] & data_operandB[20];
    assign w_20_23 = data_operandA[3] & data_operandB[20];
    assign w_20_24 = data_operandA[4] & data_operandB[20];
    assign w_20_25 = data_operandA[5] & data_operandB[20];
    assign w_20_26 = data_operandA[6] & data_operandB[20];
    assign w_20_27 = data_operandA[7] & data_operandB[20];
    assign w_20_28 = data_operandA[8] & data_operandB[20];
    assign w_20_29 = data_operandA[9] & data_operandB[20];
    assign w_20_30 = data_operandA[10] & data_operandB[20];
    assign w_20_31 = data_operandA[11] & data_operandB[20];
    assign w_20_32 = data_operandA[12] & data_operandB[20];
    assign w_20_33 = data_operandA[13] & data_operandB[20];
    assign w_20_34 = data_operandA[14] & data_operandB[20];
    assign w_20_35 = data_operandA[15] & data_operandB[20];
    assign w_20_36 = data_operandA[16] & data_operandB[20];
    assign w_20_37 = data_operandA[17] & data_operandB[20];
    assign w_20_38 = data_operandA[18] & data_operandB[20];
    assign w_20_39 = data_operandA[19] & data_operandB[20];
    assign w_20_40 = data_operandA[20] & data_operandB[20];
    assign w_20_41 = data_operandA[21] & data_operandB[20];
    assign w_20_42 = data_operandA[22] & data_operandB[20];
    assign w_20_43 = data_operandA[23] & data_operandB[20];
    assign w_20_44 = data_operandA[24] & data_operandB[20];
    assign w_20_45 = data_operandA[25] & data_operandB[20];
    assign w_20_46 = data_operandA[26] & data_operandB[20];
    assign w_20_47 = data_operandA[27] & data_operandB[20];
    assign w_20_48 = data_operandA[28] & data_operandB[20];
    assign w_20_49 = data_operandA[29] & data_operandB[20];
    assign w_20_50 = data_operandA[30] & data_operandB[20];
    assign w_20_51 = ~(data_operandA[31] & data_operandB[20]);
    full_adder adder_20_20(.S(s_20_20), .Cout(c_20_20), .A(s_19_20), .B(w_20_20), .Cin(1'b0));
    full_adder adder_20_21(.S(s_20_21), .Cout(c_20_21), .A(s_19_21), .B(w_20_21), .Cin(c_20_20));
    full_adder adder_20_22(.S(s_20_22), .Cout(c_20_22), .A(s_19_22), .B(w_20_22), .Cin(c_20_21));
    full_adder adder_20_23(.S(s_20_23), .Cout(c_20_23), .A(s_19_23), .B(w_20_23), .Cin(c_20_22));
    full_adder adder_20_24(.S(s_20_24), .Cout(c_20_24), .A(s_19_24), .B(w_20_24), .Cin(c_20_23));
    full_adder adder_20_25(.S(s_20_25), .Cout(c_20_25), .A(s_19_25), .B(w_20_25), .Cin(c_20_24));
    full_adder adder_20_26(.S(s_20_26), .Cout(c_20_26), .A(s_19_26), .B(w_20_26), .Cin(c_20_25));
    full_adder adder_20_27(.S(s_20_27), .Cout(c_20_27), .A(s_19_27), .B(w_20_27), .Cin(c_20_26));
    full_adder adder_20_28(.S(s_20_28), .Cout(c_20_28), .A(s_19_28), .B(w_20_28), .Cin(c_20_27));
    full_adder adder_20_29(.S(s_20_29), .Cout(c_20_29), .A(s_19_29), .B(w_20_29), .Cin(c_20_28));
    full_adder adder_20_30(.S(s_20_30), .Cout(c_20_30), .A(s_19_30), .B(w_20_30), .Cin(c_20_29));
    full_adder adder_20_31(.S(s_20_31), .Cout(c_20_31), .A(s_19_31), .B(w_20_31), .Cin(c_20_30));
    full_adder adder_20_32(.S(s_20_32), .Cout(c_20_32), .A(s_19_32), .B(w_20_32), .Cin(c_20_31));
    full_adder adder_20_33(.S(s_20_33), .Cout(c_20_33), .A(s_19_33), .B(w_20_33), .Cin(c_20_32));
    full_adder adder_20_34(.S(s_20_34), .Cout(c_20_34), .A(s_19_34), .B(w_20_34), .Cin(c_20_33));
    full_adder adder_20_35(.S(s_20_35), .Cout(c_20_35), .A(s_19_35), .B(w_20_35), .Cin(c_20_34));
    full_adder adder_20_36(.S(s_20_36), .Cout(c_20_36), .A(s_19_36), .B(w_20_36), .Cin(c_20_35));
    full_adder adder_20_37(.S(s_20_37), .Cout(c_20_37), .A(s_19_37), .B(w_20_37), .Cin(c_20_36));
    full_adder adder_20_38(.S(s_20_38), .Cout(c_20_38), .A(s_19_38), .B(w_20_38), .Cin(c_20_37));
    full_adder adder_20_39(.S(s_20_39), .Cout(c_20_39), .A(s_19_39), .B(w_20_39), .Cin(c_20_38));
    full_adder adder_20_40(.S(s_20_40), .Cout(c_20_40), .A(s_19_40), .B(w_20_40), .Cin(c_20_39));
    full_adder adder_20_41(.S(s_20_41), .Cout(c_20_41), .A(s_19_41), .B(w_20_41), .Cin(c_20_40));
    full_adder adder_20_42(.S(s_20_42), .Cout(c_20_42), .A(s_19_42), .B(w_20_42), .Cin(c_20_41));
    full_adder adder_20_43(.S(s_20_43), .Cout(c_20_43), .A(s_19_43), .B(w_20_43), .Cin(c_20_42));
    full_adder adder_20_44(.S(s_20_44), .Cout(c_20_44), .A(s_19_44), .B(w_20_44), .Cin(c_20_43));
    full_adder adder_20_45(.S(s_20_45), .Cout(c_20_45), .A(s_19_45), .B(w_20_45), .Cin(c_20_44));
    full_adder adder_20_46(.S(s_20_46), .Cout(c_20_46), .A(s_19_46), .B(w_20_46), .Cin(c_20_45));
    full_adder adder_20_47(.S(s_20_47), .Cout(c_20_47), .A(s_19_47), .B(w_20_47), .Cin(c_20_46));
    full_adder adder_20_48(.S(s_20_48), .Cout(c_20_48), .A(s_19_48), .B(w_20_48), .Cin(c_20_47));
    full_adder adder_20_49(.S(s_20_49), .Cout(c_20_49), .A(s_19_49), .B(w_20_49), .Cin(c_20_48));
    full_adder adder_20_50(.S(s_20_50), .Cout(c_20_50), .A(s_19_50), .B(w_20_50), .Cin(c_20_49));
    full_adder adder_20_51(.S(s_20_51), .Cout(c_20_51), .A(c_19_50), .B(w_20_51), .Cin(c_20_50));
    assign result[20] = s_20_20;
    wire w_21_21, w_21_22, w_21_23, w_21_24, w_21_25, w_21_26, w_21_27, w_21_28, w_21_29, w_21_30, w_21_31, w_21_32, w_21_33, w_21_34, w_21_35, w_21_36, w_21_37, w_21_38, w_21_39, w_21_40, w_21_41, w_21_42, w_21_43, w_21_44, w_21_45, w_21_46, w_21_47, w_21_48, w_21_49, w_21_50, w_21_51, w_21_52;
    wire s_21_21, s_21_22, s_21_23, s_21_24, s_21_25, s_21_26, s_21_27, s_21_28, s_21_29, s_21_30, s_21_31, s_21_32, s_21_33, s_21_34, s_21_35, s_21_36, s_21_37, s_21_38, s_21_39, s_21_40, s_21_41, s_21_42, s_21_43, s_21_44, s_21_45, s_21_46, s_21_47, s_21_48, s_21_49, s_21_50, s_21_51, s_21_52;
    wire c_21_21, c_21_22, c_21_23, c_21_24, c_21_25, c_21_26, c_21_27, c_21_28, c_21_29, c_21_30, c_21_31, c_21_32, c_21_33, c_21_34, c_21_35, c_21_36, c_21_37, c_21_38, c_21_39, c_21_40, c_21_41, c_21_42, c_21_43, c_21_44, c_21_45, c_21_46, c_21_47, c_21_48, c_21_49, c_21_50, c_21_51, c_21_52;
    assign w_21_21 = data_operandA[0] & data_operandB[21];
    assign w_21_22 = data_operandA[1] & data_operandB[21];
    assign w_21_23 = data_operandA[2] & data_operandB[21];
    assign w_21_24 = data_operandA[3] & data_operandB[21];
    assign w_21_25 = data_operandA[4] & data_operandB[21];
    assign w_21_26 = data_operandA[5] & data_operandB[21];
    assign w_21_27 = data_operandA[6] & data_operandB[21];
    assign w_21_28 = data_operandA[7] & data_operandB[21];
    assign w_21_29 = data_operandA[8] & data_operandB[21];
    assign w_21_30 = data_operandA[9] & data_operandB[21];
    assign w_21_31 = data_operandA[10] & data_operandB[21];
    assign w_21_32 = data_operandA[11] & data_operandB[21];
    assign w_21_33 = data_operandA[12] & data_operandB[21];
    assign w_21_34 = data_operandA[13] & data_operandB[21];
    assign w_21_35 = data_operandA[14] & data_operandB[21];
    assign w_21_36 = data_operandA[15] & data_operandB[21];
    assign w_21_37 = data_operandA[16] & data_operandB[21];
    assign w_21_38 = data_operandA[17] & data_operandB[21];
    assign w_21_39 = data_operandA[18] & data_operandB[21];
    assign w_21_40 = data_operandA[19] & data_operandB[21];
    assign w_21_41 = data_operandA[20] & data_operandB[21];
    assign w_21_42 = data_operandA[21] & data_operandB[21];
    assign w_21_43 = data_operandA[22] & data_operandB[21];
    assign w_21_44 = data_operandA[23] & data_operandB[21];
    assign w_21_45 = data_operandA[24] & data_operandB[21];
    assign w_21_46 = data_operandA[25] & data_operandB[21];
    assign w_21_47 = data_operandA[26] & data_operandB[21];
    assign w_21_48 = data_operandA[27] & data_operandB[21];
    assign w_21_49 = data_operandA[28] & data_operandB[21];
    assign w_21_50 = data_operandA[29] & data_operandB[21];
    assign w_21_51 = data_operandA[30] & data_operandB[21];
    assign w_21_52 = ~(data_operandA[31] & data_operandB[21]);
    full_adder adder_21_21(.S(s_21_21), .Cout(c_21_21), .A(s_20_21), .B(w_21_21), .Cin(1'b0));
    full_adder adder_21_22(.S(s_21_22), .Cout(c_21_22), .A(s_20_22), .B(w_21_22), .Cin(c_21_21));
    full_adder adder_21_23(.S(s_21_23), .Cout(c_21_23), .A(s_20_23), .B(w_21_23), .Cin(c_21_22));
    full_adder adder_21_24(.S(s_21_24), .Cout(c_21_24), .A(s_20_24), .B(w_21_24), .Cin(c_21_23));
    full_adder adder_21_25(.S(s_21_25), .Cout(c_21_25), .A(s_20_25), .B(w_21_25), .Cin(c_21_24));
    full_adder adder_21_26(.S(s_21_26), .Cout(c_21_26), .A(s_20_26), .B(w_21_26), .Cin(c_21_25));
    full_adder adder_21_27(.S(s_21_27), .Cout(c_21_27), .A(s_20_27), .B(w_21_27), .Cin(c_21_26));
    full_adder adder_21_28(.S(s_21_28), .Cout(c_21_28), .A(s_20_28), .B(w_21_28), .Cin(c_21_27));
    full_adder adder_21_29(.S(s_21_29), .Cout(c_21_29), .A(s_20_29), .B(w_21_29), .Cin(c_21_28));
    full_adder adder_21_30(.S(s_21_30), .Cout(c_21_30), .A(s_20_30), .B(w_21_30), .Cin(c_21_29));
    full_adder adder_21_31(.S(s_21_31), .Cout(c_21_31), .A(s_20_31), .B(w_21_31), .Cin(c_21_30));
    full_adder adder_21_32(.S(s_21_32), .Cout(c_21_32), .A(s_20_32), .B(w_21_32), .Cin(c_21_31));
    full_adder adder_21_33(.S(s_21_33), .Cout(c_21_33), .A(s_20_33), .B(w_21_33), .Cin(c_21_32));
    full_adder adder_21_34(.S(s_21_34), .Cout(c_21_34), .A(s_20_34), .B(w_21_34), .Cin(c_21_33));
    full_adder adder_21_35(.S(s_21_35), .Cout(c_21_35), .A(s_20_35), .B(w_21_35), .Cin(c_21_34));
    full_adder adder_21_36(.S(s_21_36), .Cout(c_21_36), .A(s_20_36), .B(w_21_36), .Cin(c_21_35));
    full_adder adder_21_37(.S(s_21_37), .Cout(c_21_37), .A(s_20_37), .B(w_21_37), .Cin(c_21_36));
    full_adder adder_21_38(.S(s_21_38), .Cout(c_21_38), .A(s_20_38), .B(w_21_38), .Cin(c_21_37));
    full_adder adder_21_39(.S(s_21_39), .Cout(c_21_39), .A(s_20_39), .B(w_21_39), .Cin(c_21_38));
    full_adder adder_21_40(.S(s_21_40), .Cout(c_21_40), .A(s_20_40), .B(w_21_40), .Cin(c_21_39));
    full_adder adder_21_41(.S(s_21_41), .Cout(c_21_41), .A(s_20_41), .B(w_21_41), .Cin(c_21_40));
    full_adder adder_21_42(.S(s_21_42), .Cout(c_21_42), .A(s_20_42), .B(w_21_42), .Cin(c_21_41));
    full_adder adder_21_43(.S(s_21_43), .Cout(c_21_43), .A(s_20_43), .B(w_21_43), .Cin(c_21_42));
    full_adder adder_21_44(.S(s_21_44), .Cout(c_21_44), .A(s_20_44), .B(w_21_44), .Cin(c_21_43));
    full_adder adder_21_45(.S(s_21_45), .Cout(c_21_45), .A(s_20_45), .B(w_21_45), .Cin(c_21_44));
    full_adder adder_21_46(.S(s_21_46), .Cout(c_21_46), .A(s_20_46), .B(w_21_46), .Cin(c_21_45));
    full_adder adder_21_47(.S(s_21_47), .Cout(c_21_47), .A(s_20_47), .B(w_21_47), .Cin(c_21_46));
    full_adder adder_21_48(.S(s_21_48), .Cout(c_21_48), .A(s_20_48), .B(w_21_48), .Cin(c_21_47));
    full_adder adder_21_49(.S(s_21_49), .Cout(c_21_49), .A(s_20_49), .B(w_21_49), .Cin(c_21_48));
    full_adder adder_21_50(.S(s_21_50), .Cout(c_21_50), .A(s_20_50), .B(w_21_50), .Cin(c_21_49));
    full_adder adder_21_51(.S(s_21_51), .Cout(c_21_51), .A(s_20_51), .B(w_21_51), .Cin(c_21_50));
    full_adder adder_21_52(.S(s_21_52), .Cout(c_21_52), .A(c_20_51), .B(w_21_52), .Cin(c_21_51));
    assign result[21] = s_21_21;
    wire w_22_22, w_22_23, w_22_24, w_22_25, w_22_26, w_22_27, w_22_28, w_22_29, w_22_30, w_22_31, w_22_32, w_22_33, w_22_34, w_22_35, w_22_36, w_22_37, w_22_38, w_22_39, w_22_40, w_22_41, w_22_42, w_22_43, w_22_44, w_22_45, w_22_46, w_22_47, w_22_48, w_22_49, w_22_50, w_22_51, w_22_52, w_22_53;
    wire s_22_22, s_22_23, s_22_24, s_22_25, s_22_26, s_22_27, s_22_28, s_22_29, s_22_30, s_22_31, s_22_32, s_22_33, s_22_34, s_22_35, s_22_36, s_22_37, s_22_38, s_22_39, s_22_40, s_22_41, s_22_42, s_22_43, s_22_44, s_22_45, s_22_46, s_22_47, s_22_48, s_22_49, s_22_50, s_22_51, s_22_52, s_22_53;
    wire c_22_22, c_22_23, c_22_24, c_22_25, c_22_26, c_22_27, c_22_28, c_22_29, c_22_30, c_22_31, c_22_32, c_22_33, c_22_34, c_22_35, c_22_36, c_22_37, c_22_38, c_22_39, c_22_40, c_22_41, c_22_42, c_22_43, c_22_44, c_22_45, c_22_46, c_22_47, c_22_48, c_22_49, c_22_50, c_22_51, c_22_52, c_22_53;
    assign w_22_22 = data_operandA[0] & data_operandB[22];
    assign w_22_23 = data_operandA[1] & data_operandB[22];
    assign w_22_24 = data_operandA[2] & data_operandB[22];
    assign w_22_25 = data_operandA[3] & data_operandB[22];
    assign w_22_26 = data_operandA[4] & data_operandB[22];
    assign w_22_27 = data_operandA[5] & data_operandB[22];
    assign w_22_28 = data_operandA[6] & data_operandB[22];
    assign w_22_29 = data_operandA[7] & data_operandB[22];
    assign w_22_30 = data_operandA[8] & data_operandB[22];
    assign w_22_31 = data_operandA[9] & data_operandB[22];
    assign w_22_32 = data_operandA[10] & data_operandB[22];
    assign w_22_33 = data_operandA[11] & data_operandB[22];
    assign w_22_34 = data_operandA[12] & data_operandB[22];
    assign w_22_35 = data_operandA[13] & data_operandB[22];
    assign w_22_36 = data_operandA[14] & data_operandB[22];
    assign w_22_37 = data_operandA[15] & data_operandB[22];
    assign w_22_38 = data_operandA[16] & data_operandB[22];
    assign w_22_39 = data_operandA[17] & data_operandB[22];
    assign w_22_40 = data_operandA[18] & data_operandB[22];
    assign w_22_41 = data_operandA[19] & data_operandB[22];
    assign w_22_42 = data_operandA[20] & data_operandB[22];
    assign w_22_43 = data_operandA[21] & data_operandB[22];
    assign w_22_44 = data_operandA[22] & data_operandB[22];
    assign w_22_45 = data_operandA[23] & data_operandB[22];
    assign w_22_46 = data_operandA[24] & data_operandB[22];
    assign w_22_47 = data_operandA[25] & data_operandB[22];
    assign w_22_48 = data_operandA[26] & data_operandB[22];
    assign w_22_49 = data_operandA[27] & data_operandB[22];
    assign w_22_50 = data_operandA[28] & data_operandB[22];
    assign w_22_51 = data_operandA[29] & data_operandB[22];
    assign w_22_52 = data_operandA[30] & data_operandB[22];
    assign w_22_53 = ~(data_operandA[31] & data_operandB[22]);
    full_adder adder_22_22(.S(s_22_22), .Cout(c_22_22), .A(s_21_22), .B(w_22_22), .Cin(1'b0));
    full_adder adder_22_23(.S(s_22_23), .Cout(c_22_23), .A(s_21_23), .B(w_22_23), .Cin(c_22_22));
    full_adder adder_22_24(.S(s_22_24), .Cout(c_22_24), .A(s_21_24), .B(w_22_24), .Cin(c_22_23));
    full_adder adder_22_25(.S(s_22_25), .Cout(c_22_25), .A(s_21_25), .B(w_22_25), .Cin(c_22_24));
    full_adder adder_22_26(.S(s_22_26), .Cout(c_22_26), .A(s_21_26), .B(w_22_26), .Cin(c_22_25));
    full_adder adder_22_27(.S(s_22_27), .Cout(c_22_27), .A(s_21_27), .B(w_22_27), .Cin(c_22_26));
    full_adder adder_22_28(.S(s_22_28), .Cout(c_22_28), .A(s_21_28), .B(w_22_28), .Cin(c_22_27));
    full_adder adder_22_29(.S(s_22_29), .Cout(c_22_29), .A(s_21_29), .B(w_22_29), .Cin(c_22_28));
    full_adder adder_22_30(.S(s_22_30), .Cout(c_22_30), .A(s_21_30), .B(w_22_30), .Cin(c_22_29));
    full_adder adder_22_31(.S(s_22_31), .Cout(c_22_31), .A(s_21_31), .B(w_22_31), .Cin(c_22_30));
    full_adder adder_22_32(.S(s_22_32), .Cout(c_22_32), .A(s_21_32), .B(w_22_32), .Cin(c_22_31));
    full_adder adder_22_33(.S(s_22_33), .Cout(c_22_33), .A(s_21_33), .B(w_22_33), .Cin(c_22_32));
    full_adder adder_22_34(.S(s_22_34), .Cout(c_22_34), .A(s_21_34), .B(w_22_34), .Cin(c_22_33));
    full_adder adder_22_35(.S(s_22_35), .Cout(c_22_35), .A(s_21_35), .B(w_22_35), .Cin(c_22_34));
    full_adder adder_22_36(.S(s_22_36), .Cout(c_22_36), .A(s_21_36), .B(w_22_36), .Cin(c_22_35));
    full_adder adder_22_37(.S(s_22_37), .Cout(c_22_37), .A(s_21_37), .B(w_22_37), .Cin(c_22_36));
    full_adder adder_22_38(.S(s_22_38), .Cout(c_22_38), .A(s_21_38), .B(w_22_38), .Cin(c_22_37));
    full_adder adder_22_39(.S(s_22_39), .Cout(c_22_39), .A(s_21_39), .B(w_22_39), .Cin(c_22_38));
    full_adder adder_22_40(.S(s_22_40), .Cout(c_22_40), .A(s_21_40), .B(w_22_40), .Cin(c_22_39));
    full_adder adder_22_41(.S(s_22_41), .Cout(c_22_41), .A(s_21_41), .B(w_22_41), .Cin(c_22_40));
    full_adder adder_22_42(.S(s_22_42), .Cout(c_22_42), .A(s_21_42), .B(w_22_42), .Cin(c_22_41));
    full_adder adder_22_43(.S(s_22_43), .Cout(c_22_43), .A(s_21_43), .B(w_22_43), .Cin(c_22_42));
    full_adder adder_22_44(.S(s_22_44), .Cout(c_22_44), .A(s_21_44), .B(w_22_44), .Cin(c_22_43));
    full_adder adder_22_45(.S(s_22_45), .Cout(c_22_45), .A(s_21_45), .B(w_22_45), .Cin(c_22_44));
    full_adder adder_22_46(.S(s_22_46), .Cout(c_22_46), .A(s_21_46), .B(w_22_46), .Cin(c_22_45));
    full_adder adder_22_47(.S(s_22_47), .Cout(c_22_47), .A(s_21_47), .B(w_22_47), .Cin(c_22_46));
    full_adder adder_22_48(.S(s_22_48), .Cout(c_22_48), .A(s_21_48), .B(w_22_48), .Cin(c_22_47));
    full_adder adder_22_49(.S(s_22_49), .Cout(c_22_49), .A(s_21_49), .B(w_22_49), .Cin(c_22_48));
    full_adder adder_22_50(.S(s_22_50), .Cout(c_22_50), .A(s_21_50), .B(w_22_50), .Cin(c_22_49));
    full_adder adder_22_51(.S(s_22_51), .Cout(c_22_51), .A(s_21_51), .B(w_22_51), .Cin(c_22_50));
    full_adder adder_22_52(.S(s_22_52), .Cout(c_22_52), .A(s_21_52), .B(w_22_52), .Cin(c_22_51));
    full_adder adder_22_53(.S(s_22_53), .Cout(c_22_53), .A(c_21_52), .B(w_22_53), .Cin(c_22_52));
    assign result[22] = s_22_22;
    wire w_23_23, w_23_24, w_23_25, w_23_26, w_23_27, w_23_28, w_23_29, w_23_30, w_23_31, w_23_32, w_23_33, w_23_34, w_23_35, w_23_36, w_23_37, w_23_38, w_23_39, w_23_40, w_23_41, w_23_42, w_23_43, w_23_44, w_23_45, w_23_46, w_23_47, w_23_48, w_23_49, w_23_50, w_23_51, w_23_52, w_23_53, w_23_54;
    wire s_23_23, s_23_24, s_23_25, s_23_26, s_23_27, s_23_28, s_23_29, s_23_30, s_23_31, s_23_32, s_23_33, s_23_34, s_23_35, s_23_36, s_23_37, s_23_38, s_23_39, s_23_40, s_23_41, s_23_42, s_23_43, s_23_44, s_23_45, s_23_46, s_23_47, s_23_48, s_23_49, s_23_50, s_23_51, s_23_52, s_23_53, s_23_54;
    wire c_23_23, c_23_24, c_23_25, c_23_26, c_23_27, c_23_28, c_23_29, c_23_30, c_23_31, c_23_32, c_23_33, c_23_34, c_23_35, c_23_36, c_23_37, c_23_38, c_23_39, c_23_40, c_23_41, c_23_42, c_23_43, c_23_44, c_23_45, c_23_46, c_23_47, c_23_48, c_23_49, c_23_50, c_23_51, c_23_52, c_23_53, c_23_54;
    assign w_23_23 = data_operandA[0] & data_operandB[23];
    assign w_23_24 = data_operandA[1] & data_operandB[23];
    assign w_23_25 = data_operandA[2] & data_operandB[23];
    assign w_23_26 = data_operandA[3] & data_operandB[23];
    assign w_23_27 = data_operandA[4] & data_operandB[23];
    assign w_23_28 = data_operandA[5] & data_operandB[23];
    assign w_23_29 = data_operandA[6] & data_operandB[23];
    assign w_23_30 = data_operandA[7] & data_operandB[23];
    assign w_23_31 = data_operandA[8] & data_operandB[23];
    assign w_23_32 = data_operandA[9] & data_operandB[23];
    assign w_23_33 = data_operandA[10] & data_operandB[23];
    assign w_23_34 = data_operandA[11] & data_operandB[23];
    assign w_23_35 = data_operandA[12] & data_operandB[23];
    assign w_23_36 = data_operandA[13] & data_operandB[23];
    assign w_23_37 = data_operandA[14] & data_operandB[23];
    assign w_23_38 = data_operandA[15] & data_operandB[23];
    assign w_23_39 = data_operandA[16] & data_operandB[23];
    assign w_23_40 = data_operandA[17] & data_operandB[23];
    assign w_23_41 = data_operandA[18] & data_operandB[23];
    assign w_23_42 = data_operandA[19] & data_operandB[23];
    assign w_23_43 = data_operandA[20] & data_operandB[23];
    assign w_23_44 = data_operandA[21] & data_operandB[23];
    assign w_23_45 = data_operandA[22] & data_operandB[23];
    assign w_23_46 = data_operandA[23] & data_operandB[23];
    assign w_23_47 = data_operandA[24] & data_operandB[23];
    assign w_23_48 = data_operandA[25] & data_operandB[23];
    assign w_23_49 = data_operandA[26] & data_operandB[23];
    assign w_23_50 = data_operandA[27] & data_operandB[23];
    assign w_23_51 = data_operandA[28] & data_operandB[23];
    assign w_23_52 = data_operandA[29] & data_operandB[23];
    assign w_23_53 = data_operandA[30] & data_operandB[23];
    assign w_23_54 = ~(data_operandA[31] & data_operandB[23]);
    full_adder adder_23_23(.S(s_23_23), .Cout(c_23_23), .A(s_22_23), .B(w_23_23), .Cin(1'b0));
    full_adder adder_23_24(.S(s_23_24), .Cout(c_23_24), .A(s_22_24), .B(w_23_24), .Cin(c_23_23));
    full_adder adder_23_25(.S(s_23_25), .Cout(c_23_25), .A(s_22_25), .B(w_23_25), .Cin(c_23_24));
    full_adder adder_23_26(.S(s_23_26), .Cout(c_23_26), .A(s_22_26), .B(w_23_26), .Cin(c_23_25));
    full_adder adder_23_27(.S(s_23_27), .Cout(c_23_27), .A(s_22_27), .B(w_23_27), .Cin(c_23_26));
    full_adder adder_23_28(.S(s_23_28), .Cout(c_23_28), .A(s_22_28), .B(w_23_28), .Cin(c_23_27));
    full_adder adder_23_29(.S(s_23_29), .Cout(c_23_29), .A(s_22_29), .B(w_23_29), .Cin(c_23_28));
    full_adder adder_23_30(.S(s_23_30), .Cout(c_23_30), .A(s_22_30), .B(w_23_30), .Cin(c_23_29));
    full_adder adder_23_31(.S(s_23_31), .Cout(c_23_31), .A(s_22_31), .B(w_23_31), .Cin(c_23_30));
    full_adder adder_23_32(.S(s_23_32), .Cout(c_23_32), .A(s_22_32), .B(w_23_32), .Cin(c_23_31));
    full_adder adder_23_33(.S(s_23_33), .Cout(c_23_33), .A(s_22_33), .B(w_23_33), .Cin(c_23_32));
    full_adder adder_23_34(.S(s_23_34), .Cout(c_23_34), .A(s_22_34), .B(w_23_34), .Cin(c_23_33));
    full_adder adder_23_35(.S(s_23_35), .Cout(c_23_35), .A(s_22_35), .B(w_23_35), .Cin(c_23_34));
    full_adder adder_23_36(.S(s_23_36), .Cout(c_23_36), .A(s_22_36), .B(w_23_36), .Cin(c_23_35));
    full_adder adder_23_37(.S(s_23_37), .Cout(c_23_37), .A(s_22_37), .B(w_23_37), .Cin(c_23_36));
    full_adder adder_23_38(.S(s_23_38), .Cout(c_23_38), .A(s_22_38), .B(w_23_38), .Cin(c_23_37));
    full_adder adder_23_39(.S(s_23_39), .Cout(c_23_39), .A(s_22_39), .B(w_23_39), .Cin(c_23_38));
    full_adder adder_23_40(.S(s_23_40), .Cout(c_23_40), .A(s_22_40), .B(w_23_40), .Cin(c_23_39));
    full_adder adder_23_41(.S(s_23_41), .Cout(c_23_41), .A(s_22_41), .B(w_23_41), .Cin(c_23_40));
    full_adder adder_23_42(.S(s_23_42), .Cout(c_23_42), .A(s_22_42), .B(w_23_42), .Cin(c_23_41));
    full_adder adder_23_43(.S(s_23_43), .Cout(c_23_43), .A(s_22_43), .B(w_23_43), .Cin(c_23_42));
    full_adder adder_23_44(.S(s_23_44), .Cout(c_23_44), .A(s_22_44), .B(w_23_44), .Cin(c_23_43));
    full_adder adder_23_45(.S(s_23_45), .Cout(c_23_45), .A(s_22_45), .B(w_23_45), .Cin(c_23_44));
    full_adder adder_23_46(.S(s_23_46), .Cout(c_23_46), .A(s_22_46), .B(w_23_46), .Cin(c_23_45));
    full_adder adder_23_47(.S(s_23_47), .Cout(c_23_47), .A(s_22_47), .B(w_23_47), .Cin(c_23_46));
    full_adder adder_23_48(.S(s_23_48), .Cout(c_23_48), .A(s_22_48), .B(w_23_48), .Cin(c_23_47));
    full_adder adder_23_49(.S(s_23_49), .Cout(c_23_49), .A(s_22_49), .B(w_23_49), .Cin(c_23_48));
    full_adder adder_23_50(.S(s_23_50), .Cout(c_23_50), .A(s_22_50), .B(w_23_50), .Cin(c_23_49));
    full_adder adder_23_51(.S(s_23_51), .Cout(c_23_51), .A(s_22_51), .B(w_23_51), .Cin(c_23_50));
    full_adder adder_23_52(.S(s_23_52), .Cout(c_23_52), .A(s_22_52), .B(w_23_52), .Cin(c_23_51));
    full_adder adder_23_53(.S(s_23_53), .Cout(c_23_53), .A(s_22_53), .B(w_23_53), .Cin(c_23_52));
    full_adder adder_23_54(.S(s_23_54), .Cout(c_23_54), .A(c_22_53), .B(w_23_54), .Cin(c_23_53));
    assign result[23] = s_23_23;
    wire w_24_24, w_24_25, w_24_26, w_24_27, w_24_28, w_24_29, w_24_30, w_24_31, w_24_32, w_24_33, w_24_34, w_24_35, w_24_36, w_24_37, w_24_38, w_24_39, w_24_40, w_24_41, w_24_42, w_24_43, w_24_44, w_24_45, w_24_46, w_24_47, w_24_48, w_24_49, w_24_50, w_24_51, w_24_52, w_24_53, w_24_54, w_24_55;
    wire s_24_24, s_24_25, s_24_26, s_24_27, s_24_28, s_24_29, s_24_30, s_24_31, s_24_32, s_24_33, s_24_34, s_24_35, s_24_36, s_24_37, s_24_38, s_24_39, s_24_40, s_24_41, s_24_42, s_24_43, s_24_44, s_24_45, s_24_46, s_24_47, s_24_48, s_24_49, s_24_50, s_24_51, s_24_52, s_24_53, s_24_54, s_24_55;
    wire c_24_24, c_24_25, c_24_26, c_24_27, c_24_28, c_24_29, c_24_30, c_24_31, c_24_32, c_24_33, c_24_34, c_24_35, c_24_36, c_24_37, c_24_38, c_24_39, c_24_40, c_24_41, c_24_42, c_24_43, c_24_44, c_24_45, c_24_46, c_24_47, c_24_48, c_24_49, c_24_50, c_24_51, c_24_52, c_24_53, c_24_54, c_24_55;
    assign w_24_24 = data_operandA[0] & data_operandB[24];
    assign w_24_25 = data_operandA[1] & data_operandB[24];
    assign w_24_26 = data_operandA[2] & data_operandB[24];
    assign w_24_27 = data_operandA[3] & data_operandB[24];
    assign w_24_28 = data_operandA[4] & data_operandB[24];
    assign w_24_29 = data_operandA[5] & data_operandB[24];
    assign w_24_30 = data_operandA[6] & data_operandB[24];
    assign w_24_31 = data_operandA[7] & data_operandB[24];
    assign w_24_32 = data_operandA[8] & data_operandB[24];
    assign w_24_33 = data_operandA[9] & data_operandB[24];
    assign w_24_34 = data_operandA[10] & data_operandB[24];
    assign w_24_35 = data_operandA[11] & data_operandB[24];
    assign w_24_36 = data_operandA[12] & data_operandB[24];
    assign w_24_37 = data_operandA[13] & data_operandB[24];
    assign w_24_38 = data_operandA[14] & data_operandB[24];
    assign w_24_39 = data_operandA[15] & data_operandB[24];
    assign w_24_40 = data_operandA[16] & data_operandB[24];
    assign w_24_41 = data_operandA[17] & data_operandB[24];
    assign w_24_42 = data_operandA[18] & data_operandB[24];
    assign w_24_43 = data_operandA[19] & data_operandB[24];
    assign w_24_44 = data_operandA[20] & data_operandB[24];
    assign w_24_45 = data_operandA[21] & data_operandB[24];
    assign w_24_46 = data_operandA[22] & data_operandB[24];
    assign w_24_47 = data_operandA[23] & data_operandB[24];
    assign w_24_48 = data_operandA[24] & data_operandB[24];
    assign w_24_49 = data_operandA[25] & data_operandB[24];
    assign w_24_50 = data_operandA[26] & data_operandB[24];
    assign w_24_51 = data_operandA[27] & data_operandB[24];
    assign w_24_52 = data_operandA[28] & data_operandB[24];
    assign w_24_53 = data_operandA[29] & data_operandB[24];
    assign w_24_54 = data_operandA[30] & data_operandB[24];
    assign w_24_55 = ~(data_operandA[31] & data_operandB[24]);
    full_adder adder_24_24(.S(s_24_24), .Cout(c_24_24), .A(s_23_24), .B(w_24_24), .Cin(1'b0));
    full_adder adder_24_25(.S(s_24_25), .Cout(c_24_25), .A(s_23_25), .B(w_24_25), .Cin(c_24_24));
    full_adder adder_24_26(.S(s_24_26), .Cout(c_24_26), .A(s_23_26), .B(w_24_26), .Cin(c_24_25));
    full_adder adder_24_27(.S(s_24_27), .Cout(c_24_27), .A(s_23_27), .B(w_24_27), .Cin(c_24_26));
    full_adder adder_24_28(.S(s_24_28), .Cout(c_24_28), .A(s_23_28), .B(w_24_28), .Cin(c_24_27));
    full_adder adder_24_29(.S(s_24_29), .Cout(c_24_29), .A(s_23_29), .B(w_24_29), .Cin(c_24_28));
    full_adder adder_24_30(.S(s_24_30), .Cout(c_24_30), .A(s_23_30), .B(w_24_30), .Cin(c_24_29));
    full_adder adder_24_31(.S(s_24_31), .Cout(c_24_31), .A(s_23_31), .B(w_24_31), .Cin(c_24_30));
    full_adder adder_24_32(.S(s_24_32), .Cout(c_24_32), .A(s_23_32), .B(w_24_32), .Cin(c_24_31));
    full_adder adder_24_33(.S(s_24_33), .Cout(c_24_33), .A(s_23_33), .B(w_24_33), .Cin(c_24_32));
    full_adder adder_24_34(.S(s_24_34), .Cout(c_24_34), .A(s_23_34), .B(w_24_34), .Cin(c_24_33));
    full_adder adder_24_35(.S(s_24_35), .Cout(c_24_35), .A(s_23_35), .B(w_24_35), .Cin(c_24_34));
    full_adder adder_24_36(.S(s_24_36), .Cout(c_24_36), .A(s_23_36), .B(w_24_36), .Cin(c_24_35));
    full_adder adder_24_37(.S(s_24_37), .Cout(c_24_37), .A(s_23_37), .B(w_24_37), .Cin(c_24_36));
    full_adder adder_24_38(.S(s_24_38), .Cout(c_24_38), .A(s_23_38), .B(w_24_38), .Cin(c_24_37));
    full_adder adder_24_39(.S(s_24_39), .Cout(c_24_39), .A(s_23_39), .B(w_24_39), .Cin(c_24_38));
    full_adder adder_24_40(.S(s_24_40), .Cout(c_24_40), .A(s_23_40), .B(w_24_40), .Cin(c_24_39));
    full_adder adder_24_41(.S(s_24_41), .Cout(c_24_41), .A(s_23_41), .B(w_24_41), .Cin(c_24_40));
    full_adder adder_24_42(.S(s_24_42), .Cout(c_24_42), .A(s_23_42), .B(w_24_42), .Cin(c_24_41));
    full_adder adder_24_43(.S(s_24_43), .Cout(c_24_43), .A(s_23_43), .B(w_24_43), .Cin(c_24_42));
    full_adder adder_24_44(.S(s_24_44), .Cout(c_24_44), .A(s_23_44), .B(w_24_44), .Cin(c_24_43));
    full_adder adder_24_45(.S(s_24_45), .Cout(c_24_45), .A(s_23_45), .B(w_24_45), .Cin(c_24_44));
    full_adder adder_24_46(.S(s_24_46), .Cout(c_24_46), .A(s_23_46), .B(w_24_46), .Cin(c_24_45));
    full_adder adder_24_47(.S(s_24_47), .Cout(c_24_47), .A(s_23_47), .B(w_24_47), .Cin(c_24_46));
    full_adder adder_24_48(.S(s_24_48), .Cout(c_24_48), .A(s_23_48), .B(w_24_48), .Cin(c_24_47));
    full_adder adder_24_49(.S(s_24_49), .Cout(c_24_49), .A(s_23_49), .B(w_24_49), .Cin(c_24_48));
    full_adder adder_24_50(.S(s_24_50), .Cout(c_24_50), .A(s_23_50), .B(w_24_50), .Cin(c_24_49));
    full_adder adder_24_51(.S(s_24_51), .Cout(c_24_51), .A(s_23_51), .B(w_24_51), .Cin(c_24_50));
    full_adder adder_24_52(.S(s_24_52), .Cout(c_24_52), .A(s_23_52), .B(w_24_52), .Cin(c_24_51));
    full_adder adder_24_53(.S(s_24_53), .Cout(c_24_53), .A(s_23_53), .B(w_24_53), .Cin(c_24_52));
    full_adder adder_24_54(.S(s_24_54), .Cout(c_24_54), .A(s_23_54), .B(w_24_54), .Cin(c_24_53));
    full_adder adder_24_55(.S(s_24_55), .Cout(c_24_55), .A(c_23_54), .B(w_24_55), .Cin(c_24_54));
    assign result[24] = s_24_24;
    wire w_25_25, w_25_26, w_25_27, w_25_28, w_25_29, w_25_30, w_25_31, w_25_32, w_25_33, w_25_34, w_25_35, w_25_36, w_25_37, w_25_38, w_25_39, w_25_40, w_25_41, w_25_42, w_25_43, w_25_44, w_25_45, w_25_46, w_25_47, w_25_48, w_25_49, w_25_50, w_25_51, w_25_52, w_25_53, w_25_54, w_25_55, w_25_56;
    wire s_25_25, s_25_26, s_25_27, s_25_28, s_25_29, s_25_30, s_25_31, s_25_32, s_25_33, s_25_34, s_25_35, s_25_36, s_25_37, s_25_38, s_25_39, s_25_40, s_25_41, s_25_42, s_25_43, s_25_44, s_25_45, s_25_46, s_25_47, s_25_48, s_25_49, s_25_50, s_25_51, s_25_52, s_25_53, s_25_54, s_25_55, s_25_56;
    wire c_25_25, c_25_26, c_25_27, c_25_28, c_25_29, c_25_30, c_25_31, c_25_32, c_25_33, c_25_34, c_25_35, c_25_36, c_25_37, c_25_38, c_25_39, c_25_40, c_25_41, c_25_42, c_25_43, c_25_44, c_25_45, c_25_46, c_25_47, c_25_48, c_25_49, c_25_50, c_25_51, c_25_52, c_25_53, c_25_54, c_25_55, c_25_56;
    assign w_25_25 = data_operandA[0] & data_operandB[25];
    assign w_25_26 = data_operandA[1] & data_operandB[25];
    assign w_25_27 = data_operandA[2] & data_operandB[25];
    assign w_25_28 = data_operandA[3] & data_operandB[25];
    assign w_25_29 = data_operandA[4] & data_operandB[25];
    assign w_25_30 = data_operandA[5] & data_operandB[25];
    assign w_25_31 = data_operandA[6] & data_operandB[25];
    assign w_25_32 = data_operandA[7] & data_operandB[25];
    assign w_25_33 = data_operandA[8] & data_operandB[25];
    assign w_25_34 = data_operandA[9] & data_operandB[25];
    assign w_25_35 = data_operandA[10] & data_operandB[25];
    assign w_25_36 = data_operandA[11] & data_operandB[25];
    assign w_25_37 = data_operandA[12] & data_operandB[25];
    assign w_25_38 = data_operandA[13] & data_operandB[25];
    assign w_25_39 = data_operandA[14] & data_operandB[25];
    assign w_25_40 = data_operandA[15] & data_operandB[25];
    assign w_25_41 = data_operandA[16] & data_operandB[25];
    assign w_25_42 = data_operandA[17] & data_operandB[25];
    assign w_25_43 = data_operandA[18] & data_operandB[25];
    assign w_25_44 = data_operandA[19] & data_operandB[25];
    assign w_25_45 = data_operandA[20] & data_operandB[25];
    assign w_25_46 = data_operandA[21] & data_operandB[25];
    assign w_25_47 = data_operandA[22] & data_operandB[25];
    assign w_25_48 = data_operandA[23] & data_operandB[25];
    assign w_25_49 = data_operandA[24] & data_operandB[25];
    assign w_25_50 = data_operandA[25] & data_operandB[25];
    assign w_25_51 = data_operandA[26] & data_operandB[25];
    assign w_25_52 = data_operandA[27] & data_operandB[25];
    assign w_25_53 = data_operandA[28] & data_operandB[25];
    assign w_25_54 = data_operandA[29] & data_operandB[25];
    assign w_25_55 = data_operandA[30] & data_operandB[25];
    assign w_25_56 = ~(data_operandA[31] & data_operandB[25]);
    full_adder adder_25_25(.S(s_25_25), .Cout(c_25_25), .A(s_24_25), .B(w_25_25), .Cin(1'b0));
    full_adder adder_25_26(.S(s_25_26), .Cout(c_25_26), .A(s_24_26), .B(w_25_26), .Cin(c_25_25));
    full_adder adder_25_27(.S(s_25_27), .Cout(c_25_27), .A(s_24_27), .B(w_25_27), .Cin(c_25_26));
    full_adder adder_25_28(.S(s_25_28), .Cout(c_25_28), .A(s_24_28), .B(w_25_28), .Cin(c_25_27));
    full_adder adder_25_29(.S(s_25_29), .Cout(c_25_29), .A(s_24_29), .B(w_25_29), .Cin(c_25_28));
    full_adder adder_25_30(.S(s_25_30), .Cout(c_25_30), .A(s_24_30), .B(w_25_30), .Cin(c_25_29));
    full_adder adder_25_31(.S(s_25_31), .Cout(c_25_31), .A(s_24_31), .B(w_25_31), .Cin(c_25_30));
    full_adder adder_25_32(.S(s_25_32), .Cout(c_25_32), .A(s_24_32), .B(w_25_32), .Cin(c_25_31));
    full_adder adder_25_33(.S(s_25_33), .Cout(c_25_33), .A(s_24_33), .B(w_25_33), .Cin(c_25_32));
    full_adder adder_25_34(.S(s_25_34), .Cout(c_25_34), .A(s_24_34), .B(w_25_34), .Cin(c_25_33));
    full_adder adder_25_35(.S(s_25_35), .Cout(c_25_35), .A(s_24_35), .B(w_25_35), .Cin(c_25_34));
    full_adder adder_25_36(.S(s_25_36), .Cout(c_25_36), .A(s_24_36), .B(w_25_36), .Cin(c_25_35));
    full_adder adder_25_37(.S(s_25_37), .Cout(c_25_37), .A(s_24_37), .B(w_25_37), .Cin(c_25_36));
    full_adder adder_25_38(.S(s_25_38), .Cout(c_25_38), .A(s_24_38), .B(w_25_38), .Cin(c_25_37));
    full_adder adder_25_39(.S(s_25_39), .Cout(c_25_39), .A(s_24_39), .B(w_25_39), .Cin(c_25_38));
    full_adder adder_25_40(.S(s_25_40), .Cout(c_25_40), .A(s_24_40), .B(w_25_40), .Cin(c_25_39));
    full_adder adder_25_41(.S(s_25_41), .Cout(c_25_41), .A(s_24_41), .B(w_25_41), .Cin(c_25_40));
    full_adder adder_25_42(.S(s_25_42), .Cout(c_25_42), .A(s_24_42), .B(w_25_42), .Cin(c_25_41));
    full_adder adder_25_43(.S(s_25_43), .Cout(c_25_43), .A(s_24_43), .B(w_25_43), .Cin(c_25_42));
    full_adder adder_25_44(.S(s_25_44), .Cout(c_25_44), .A(s_24_44), .B(w_25_44), .Cin(c_25_43));
    full_adder adder_25_45(.S(s_25_45), .Cout(c_25_45), .A(s_24_45), .B(w_25_45), .Cin(c_25_44));
    full_adder adder_25_46(.S(s_25_46), .Cout(c_25_46), .A(s_24_46), .B(w_25_46), .Cin(c_25_45));
    full_adder adder_25_47(.S(s_25_47), .Cout(c_25_47), .A(s_24_47), .B(w_25_47), .Cin(c_25_46));
    full_adder adder_25_48(.S(s_25_48), .Cout(c_25_48), .A(s_24_48), .B(w_25_48), .Cin(c_25_47));
    full_adder adder_25_49(.S(s_25_49), .Cout(c_25_49), .A(s_24_49), .B(w_25_49), .Cin(c_25_48));
    full_adder adder_25_50(.S(s_25_50), .Cout(c_25_50), .A(s_24_50), .B(w_25_50), .Cin(c_25_49));
    full_adder adder_25_51(.S(s_25_51), .Cout(c_25_51), .A(s_24_51), .B(w_25_51), .Cin(c_25_50));
    full_adder adder_25_52(.S(s_25_52), .Cout(c_25_52), .A(s_24_52), .B(w_25_52), .Cin(c_25_51));
    full_adder adder_25_53(.S(s_25_53), .Cout(c_25_53), .A(s_24_53), .B(w_25_53), .Cin(c_25_52));
    full_adder adder_25_54(.S(s_25_54), .Cout(c_25_54), .A(s_24_54), .B(w_25_54), .Cin(c_25_53));
    full_adder adder_25_55(.S(s_25_55), .Cout(c_25_55), .A(s_24_55), .B(w_25_55), .Cin(c_25_54));
    full_adder adder_25_56(.S(s_25_56), .Cout(c_25_56), .A(c_24_55), .B(w_25_56), .Cin(c_25_55));
    assign result[25] = s_25_25;
    wire w_26_26, w_26_27, w_26_28, w_26_29, w_26_30, w_26_31, w_26_32, w_26_33, w_26_34, w_26_35, w_26_36, w_26_37, w_26_38, w_26_39, w_26_40, w_26_41, w_26_42, w_26_43, w_26_44, w_26_45, w_26_46, w_26_47, w_26_48, w_26_49, w_26_50, w_26_51, w_26_52, w_26_53, w_26_54, w_26_55, w_26_56, w_26_57;
    wire s_26_26, s_26_27, s_26_28, s_26_29, s_26_30, s_26_31, s_26_32, s_26_33, s_26_34, s_26_35, s_26_36, s_26_37, s_26_38, s_26_39, s_26_40, s_26_41, s_26_42, s_26_43, s_26_44, s_26_45, s_26_46, s_26_47, s_26_48, s_26_49, s_26_50, s_26_51, s_26_52, s_26_53, s_26_54, s_26_55, s_26_56, s_26_57;
    wire c_26_26, c_26_27, c_26_28, c_26_29, c_26_30, c_26_31, c_26_32, c_26_33, c_26_34, c_26_35, c_26_36, c_26_37, c_26_38, c_26_39, c_26_40, c_26_41, c_26_42, c_26_43, c_26_44, c_26_45, c_26_46, c_26_47, c_26_48, c_26_49, c_26_50, c_26_51, c_26_52, c_26_53, c_26_54, c_26_55, c_26_56, c_26_57;
    assign w_26_26 = data_operandA[0] & data_operandB[26];
    assign w_26_27 = data_operandA[1] & data_operandB[26];
    assign w_26_28 = data_operandA[2] & data_operandB[26];
    assign w_26_29 = data_operandA[3] & data_operandB[26];
    assign w_26_30 = data_operandA[4] & data_operandB[26];
    assign w_26_31 = data_operandA[5] & data_operandB[26];
    assign w_26_32 = data_operandA[6] & data_operandB[26];
    assign w_26_33 = data_operandA[7] & data_operandB[26];
    assign w_26_34 = data_operandA[8] & data_operandB[26];
    assign w_26_35 = data_operandA[9] & data_operandB[26];
    assign w_26_36 = data_operandA[10] & data_operandB[26];
    assign w_26_37 = data_operandA[11] & data_operandB[26];
    assign w_26_38 = data_operandA[12] & data_operandB[26];
    assign w_26_39 = data_operandA[13] & data_operandB[26];
    assign w_26_40 = data_operandA[14] & data_operandB[26];
    assign w_26_41 = data_operandA[15] & data_operandB[26];
    assign w_26_42 = data_operandA[16] & data_operandB[26];
    assign w_26_43 = data_operandA[17] & data_operandB[26];
    assign w_26_44 = data_operandA[18] & data_operandB[26];
    assign w_26_45 = data_operandA[19] & data_operandB[26];
    assign w_26_46 = data_operandA[20] & data_operandB[26];
    assign w_26_47 = data_operandA[21] & data_operandB[26];
    assign w_26_48 = data_operandA[22] & data_operandB[26];
    assign w_26_49 = data_operandA[23] & data_operandB[26];
    assign w_26_50 = data_operandA[24] & data_operandB[26];
    assign w_26_51 = data_operandA[25] & data_operandB[26];
    assign w_26_52 = data_operandA[26] & data_operandB[26];
    assign w_26_53 = data_operandA[27] & data_operandB[26];
    assign w_26_54 = data_operandA[28] & data_operandB[26];
    assign w_26_55 = data_operandA[29] & data_operandB[26];
    assign w_26_56 = data_operandA[30] & data_operandB[26];
    assign w_26_57 = ~(data_operandA[31] & data_operandB[26]);
    full_adder adder_26_26(.S(s_26_26), .Cout(c_26_26), .A(s_25_26), .B(w_26_26), .Cin(1'b0));
    full_adder adder_26_27(.S(s_26_27), .Cout(c_26_27), .A(s_25_27), .B(w_26_27), .Cin(c_26_26));
    full_adder adder_26_28(.S(s_26_28), .Cout(c_26_28), .A(s_25_28), .B(w_26_28), .Cin(c_26_27));
    full_adder adder_26_29(.S(s_26_29), .Cout(c_26_29), .A(s_25_29), .B(w_26_29), .Cin(c_26_28));
    full_adder adder_26_30(.S(s_26_30), .Cout(c_26_30), .A(s_25_30), .B(w_26_30), .Cin(c_26_29));
    full_adder adder_26_31(.S(s_26_31), .Cout(c_26_31), .A(s_25_31), .B(w_26_31), .Cin(c_26_30));
    full_adder adder_26_32(.S(s_26_32), .Cout(c_26_32), .A(s_25_32), .B(w_26_32), .Cin(c_26_31));
    full_adder adder_26_33(.S(s_26_33), .Cout(c_26_33), .A(s_25_33), .B(w_26_33), .Cin(c_26_32));
    full_adder adder_26_34(.S(s_26_34), .Cout(c_26_34), .A(s_25_34), .B(w_26_34), .Cin(c_26_33));
    full_adder adder_26_35(.S(s_26_35), .Cout(c_26_35), .A(s_25_35), .B(w_26_35), .Cin(c_26_34));
    full_adder adder_26_36(.S(s_26_36), .Cout(c_26_36), .A(s_25_36), .B(w_26_36), .Cin(c_26_35));
    full_adder adder_26_37(.S(s_26_37), .Cout(c_26_37), .A(s_25_37), .B(w_26_37), .Cin(c_26_36));
    full_adder adder_26_38(.S(s_26_38), .Cout(c_26_38), .A(s_25_38), .B(w_26_38), .Cin(c_26_37));
    full_adder adder_26_39(.S(s_26_39), .Cout(c_26_39), .A(s_25_39), .B(w_26_39), .Cin(c_26_38));
    full_adder adder_26_40(.S(s_26_40), .Cout(c_26_40), .A(s_25_40), .B(w_26_40), .Cin(c_26_39));
    full_adder adder_26_41(.S(s_26_41), .Cout(c_26_41), .A(s_25_41), .B(w_26_41), .Cin(c_26_40));
    full_adder adder_26_42(.S(s_26_42), .Cout(c_26_42), .A(s_25_42), .B(w_26_42), .Cin(c_26_41));
    full_adder adder_26_43(.S(s_26_43), .Cout(c_26_43), .A(s_25_43), .B(w_26_43), .Cin(c_26_42));
    full_adder adder_26_44(.S(s_26_44), .Cout(c_26_44), .A(s_25_44), .B(w_26_44), .Cin(c_26_43));
    full_adder adder_26_45(.S(s_26_45), .Cout(c_26_45), .A(s_25_45), .B(w_26_45), .Cin(c_26_44));
    full_adder adder_26_46(.S(s_26_46), .Cout(c_26_46), .A(s_25_46), .B(w_26_46), .Cin(c_26_45));
    full_adder adder_26_47(.S(s_26_47), .Cout(c_26_47), .A(s_25_47), .B(w_26_47), .Cin(c_26_46));
    full_adder adder_26_48(.S(s_26_48), .Cout(c_26_48), .A(s_25_48), .B(w_26_48), .Cin(c_26_47));
    full_adder adder_26_49(.S(s_26_49), .Cout(c_26_49), .A(s_25_49), .B(w_26_49), .Cin(c_26_48));
    full_adder adder_26_50(.S(s_26_50), .Cout(c_26_50), .A(s_25_50), .B(w_26_50), .Cin(c_26_49));
    full_adder adder_26_51(.S(s_26_51), .Cout(c_26_51), .A(s_25_51), .B(w_26_51), .Cin(c_26_50));
    full_adder adder_26_52(.S(s_26_52), .Cout(c_26_52), .A(s_25_52), .B(w_26_52), .Cin(c_26_51));
    full_adder adder_26_53(.S(s_26_53), .Cout(c_26_53), .A(s_25_53), .B(w_26_53), .Cin(c_26_52));
    full_adder adder_26_54(.S(s_26_54), .Cout(c_26_54), .A(s_25_54), .B(w_26_54), .Cin(c_26_53));
    full_adder adder_26_55(.S(s_26_55), .Cout(c_26_55), .A(s_25_55), .B(w_26_55), .Cin(c_26_54));
    full_adder adder_26_56(.S(s_26_56), .Cout(c_26_56), .A(s_25_56), .B(w_26_56), .Cin(c_26_55));
    full_adder adder_26_57(.S(s_26_57), .Cout(c_26_57), .A(c_25_56), .B(w_26_57), .Cin(c_26_56));
    assign result[26] = s_26_26;
    wire w_27_27, w_27_28, w_27_29, w_27_30, w_27_31, w_27_32, w_27_33, w_27_34, w_27_35, w_27_36, w_27_37, w_27_38, w_27_39, w_27_40, w_27_41, w_27_42, w_27_43, w_27_44, w_27_45, w_27_46, w_27_47, w_27_48, w_27_49, w_27_50, w_27_51, w_27_52, w_27_53, w_27_54, w_27_55, w_27_56, w_27_57, w_27_58;
    wire s_27_27, s_27_28, s_27_29, s_27_30, s_27_31, s_27_32, s_27_33, s_27_34, s_27_35, s_27_36, s_27_37, s_27_38, s_27_39, s_27_40, s_27_41, s_27_42, s_27_43, s_27_44, s_27_45, s_27_46, s_27_47, s_27_48, s_27_49, s_27_50, s_27_51, s_27_52, s_27_53, s_27_54, s_27_55, s_27_56, s_27_57, s_27_58;
    wire c_27_27, c_27_28, c_27_29, c_27_30, c_27_31, c_27_32, c_27_33, c_27_34, c_27_35, c_27_36, c_27_37, c_27_38, c_27_39, c_27_40, c_27_41, c_27_42, c_27_43, c_27_44, c_27_45, c_27_46, c_27_47, c_27_48, c_27_49, c_27_50, c_27_51, c_27_52, c_27_53, c_27_54, c_27_55, c_27_56, c_27_57, c_27_58;
    assign w_27_27 = data_operandA[0] & data_operandB[27];
    assign w_27_28 = data_operandA[1] & data_operandB[27];
    assign w_27_29 = data_operandA[2] & data_operandB[27];
    assign w_27_30 = data_operandA[3] & data_operandB[27];
    assign w_27_31 = data_operandA[4] & data_operandB[27];
    assign w_27_32 = data_operandA[5] & data_operandB[27];
    assign w_27_33 = data_operandA[6] & data_operandB[27];
    assign w_27_34 = data_operandA[7] & data_operandB[27];
    assign w_27_35 = data_operandA[8] & data_operandB[27];
    assign w_27_36 = data_operandA[9] & data_operandB[27];
    assign w_27_37 = data_operandA[10] & data_operandB[27];
    assign w_27_38 = data_operandA[11] & data_operandB[27];
    assign w_27_39 = data_operandA[12] & data_operandB[27];
    assign w_27_40 = data_operandA[13] & data_operandB[27];
    assign w_27_41 = data_operandA[14] & data_operandB[27];
    assign w_27_42 = data_operandA[15] & data_operandB[27];
    assign w_27_43 = data_operandA[16] & data_operandB[27];
    assign w_27_44 = data_operandA[17] & data_operandB[27];
    assign w_27_45 = data_operandA[18] & data_operandB[27];
    assign w_27_46 = data_operandA[19] & data_operandB[27];
    assign w_27_47 = data_operandA[20] & data_operandB[27];
    assign w_27_48 = data_operandA[21] & data_operandB[27];
    assign w_27_49 = data_operandA[22] & data_operandB[27];
    assign w_27_50 = data_operandA[23] & data_operandB[27];
    assign w_27_51 = data_operandA[24] & data_operandB[27];
    assign w_27_52 = data_operandA[25] & data_operandB[27];
    assign w_27_53 = data_operandA[26] & data_operandB[27];
    assign w_27_54 = data_operandA[27] & data_operandB[27];
    assign w_27_55 = data_operandA[28] & data_operandB[27];
    assign w_27_56 = data_operandA[29] & data_operandB[27];
    assign w_27_57 = data_operandA[30] & data_operandB[27];
    assign w_27_58 = ~(data_operandA[31] & data_operandB[27]);
    full_adder adder_27_27(.S(s_27_27), .Cout(c_27_27), .A(s_26_27), .B(w_27_27), .Cin(1'b0));
    full_adder adder_27_28(.S(s_27_28), .Cout(c_27_28), .A(s_26_28), .B(w_27_28), .Cin(c_27_27));
    full_adder adder_27_29(.S(s_27_29), .Cout(c_27_29), .A(s_26_29), .B(w_27_29), .Cin(c_27_28));
    full_adder adder_27_30(.S(s_27_30), .Cout(c_27_30), .A(s_26_30), .B(w_27_30), .Cin(c_27_29));
    full_adder adder_27_31(.S(s_27_31), .Cout(c_27_31), .A(s_26_31), .B(w_27_31), .Cin(c_27_30));
    full_adder adder_27_32(.S(s_27_32), .Cout(c_27_32), .A(s_26_32), .B(w_27_32), .Cin(c_27_31));
    full_adder adder_27_33(.S(s_27_33), .Cout(c_27_33), .A(s_26_33), .B(w_27_33), .Cin(c_27_32));
    full_adder adder_27_34(.S(s_27_34), .Cout(c_27_34), .A(s_26_34), .B(w_27_34), .Cin(c_27_33));
    full_adder adder_27_35(.S(s_27_35), .Cout(c_27_35), .A(s_26_35), .B(w_27_35), .Cin(c_27_34));
    full_adder adder_27_36(.S(s_27_36), .Cout(c_27_36), .A(s_26_36), .B(w_27_36), .Cin(c_27_35));
    full_adder adder_27_37(.S(s_27_37), .Cout(c_27_37), .A(s_26_37), .B(w_27_37), .Cin(c_27_36));
    full_adder adder_27_38(.S(s_27_38), .Cout(c_27_38), .A(s_26_38), .B(w_27_38), .Cin(c_27_37));
    full_adder adder_27_39(.S(s_27_39), .Cout(c_27_39), .A(s_26_39), .B(w_27_39), .Cin(c_27_38));
    full_adder adder_27_40(.S(s_27_40), .Cout(c_27_40), .A(s_26_40), .B(w_27_40), .Cin(c_27_39));
    full_adder adder_27_41(.S(s_27_41), .Cout(c_27_41), .A(s_26_41), .B(w_27_41), .Cin(c_27_40));
    full_adder adder_27_42(.S(s_27_42), .Cout(c_27_42), .A(s_26_42), .B(w_27_42), .Cin(c_27_41));
    full_adder adder_27_43(.S(s_27_43), .Cout(c_27_43), .A(s_26_43), .B(w_27_43), .Cin(c_27_42));
    full_adder adder_27_44(.S(s_27_44), .Cout(c_27_44), .A(s_26_44), .B(w_27_44), .Cin(c_27_43));
    full_adder adder_27_45(.S(s_27_45), .Cout(c_27_45), .A(s_26_45), .B(w_27_45), .Cin(c_27_44));
    full_adder adder_27_46(.S(s_27_46), .Cout(c_27_46), .A(s_26_46), .B(w_27_46), .Cin(c_27_45));
    full_adder adder_27_47(.S(s_27_47), .Cout(c_27_47), .A(s_26_47), .B(w_27_47), .Cin(c_27_46));
    full_adder adder_27_48(.S(s_27_48), .Cout(c_27_48), .A(s_26_48), .B(w_27_48), .Cin(c_27_47));
    full_adder adder_27_49(.S(s_27_49), .Cout(c_27_49), .A(s_26_49), .B(w_27_49), .Cin(c_27_48));
    full_adder adder_27_50(.S(s_27_50), .Cout(c_27_50), .A(s_26_50), .B(w_27_50), .Cin(c_27_49));
    full_adder adder_27_51(.S(s_27_51), .Cout(c_27_51), .A(s_26_51), .B(w_27_51), .Cin(c_27_50));
    full_adder adder_27_52(.S(s_27_52), .Cout(c_27_52), .A(s_26_52), .B(w_27_52), .Cin(c_27_51));
    full_adder adder_27_53(.S(s_27_53), .Cout(c_27_53), .A(s_26_53), .B(w_27_53), .Cin(c_27_52));
    full_adder adder_27_54(.S(s_27_54), .Cout(c_27_54), .A(s_26_54), .B(w_27_54), .Cin(c_27_53));
    full_adder adder_27_55(.S(s_27_55), .Cout(c_27_55), .A(s_26_55), .B(w_27_55), .Cin(c_27_54));
    full_adder adder_27_56(.S(s_27_56), .Cout(c_27_56), .A(s_26_56), .B(w_27_56), .Cin(c_27_55));
    full_adder adder_27_57(.S(s_27_57), .Cout(c_27_57), .A(s_26_57), .B(w_27_57), .Cin(c_27_56));
    full_adder adder_27_58(.S(s_27_58), .Cout(c_27_58), .A(c_26_57), .B(w_27_58), .Cin(c_27_57));
    assign result[27] = s_27_27;
    wire w_28_28, w_28_29, w_28_30, w_28_31, w_28_32, w_28_33, w_28_34, w_28_35, w_28_36, w_28_37, w_28_38, w_28_39, w_28_40, w_28_41, w_28_42, w_28_43, w_28_44, w_28_45, w_28_46, w_28_47, w_28_48, w_28_49, w_28_50, w_28_51, w_28_52, w_28_53, w_28_54, w_28_55, w_28_56, w_28_57, w_28_58, w_28_59;
    wire s_28_28, s_28_29, s_28_30, s_28_31, s_28_32, s_28_33, s_28_34, s_28_35, s_28_36, s_28_37, s_28_38, s_28_39, s_28_40, s_28_41, s_28_42, s_28_43, s_28_44, s_28_45, s_28_46, s_28_47, s_28_48, s_28_49, s_28_50, s_28_51, s_28_52, s_28_53, s_28_54, s_28_55, s_28_56, s_28_57, s_28_58, s_28_59;
    wire c_28_28, c_28_29, c_28_30, c_28_31, c_28_32, c_28_33, c_28_34, c_28_35, c_28_36, c_28_37, c_28_38, c_28_39, c_28_40, c_28_41, c_28_42, c_28_43, c_28_44, c_28_45, c_28_46, c_28_47, c_28_48, c_28_49, c_28_50, c_28_51, c_28_52, c_28_53, c_28_54, c_28_55, c_28_56, c_28_57, c_28_58, c_28_59;
    assign w_28_28 = data_operandA[0] & data_operandB[28];
    assign w_28_29 = data_operandA[1] & data_operandB[28];
    assign w_28_30 = data_operandA[2] & data_operandB[28];
    assign w_28_31 = data_operandA[3] & data_operandB[28];
    assign w_28_32 = data_operandA[4] & data_operandB[28];
    assign w_28_33 = data_operandA[5] & data_operandB[28];
    assign w_28_34 = data_operandA[6] & data_operandB[28];
    assign w_28_35 = data_operandA[7] & data_operandB[28];
    assign w_28_36 = data_operandA[8] & data_operandB[28];
    assign w_28_37 = data_operandA[9] & data_operandB[28];
    assign w_28_38 = data_operandA[10] & data_operandB[28];
    assign w_28_39 = data_operandA[11] & data_operandB[28];
    assign w_28_40 = data_operandA[12] & data_operandB[28];
    assign w_28_41 = data_operandA[13] & data_operandB[28];
    assign w_28_42 = data_operandA[14] & data_operandB[28];
    assign w_28_43 = data_operandA[15] & data_operandB[28];
    assign w_28_44 = data_operandA[16] & data_operandB[28];
    assign w_28_45 = data_operandA[17] & data_operandB[28];
    assign w_28_46 = data_operandA[18] & data_operandB[28];
    assign w_28_47 = data_operandA[19] & data_operandB[28];
    assign w_28_48 = data_operandA[20] & data_operandB[28];
    assign w_28_49 = data_operandA[21] & data_operandB[28];
    assign w_28_50 = data_operandA[22] & data_operandB[28];
    assign w_28_51 = data_operandA[23] & data_operandB[28];
    assign w_28_52 = data_operandA[24] & data_operandB[28];
    assign w_28_53 = data_operandA[25] & data_operandB[28];
    assign w_28_54 = data_operandA[26] & data_operandB[28];
    assign w_28_55 = data_operandA[27] & data_operandB[28];
    assign w_28_56 = data_operandA[28] & data_operandB[28];
    assign w_28_57 = data_operandA[29] & data_operandB[28];
    assign w_28_58 = data_operandA[30] & data_operandB[28];
    assign w_28_59 = ~(data_operandA[31] & data_operandB[28]);
    full_adder adder_28_28(.S(s_28_28), .Cout(c_28_28), .A(s_27_28), .B(w_28_28), .Cin(1'b0));
    full_adder adder_28_29(.S(s_28_29), .Cout(c_28_29), .A(s_27_29), .B(w_28_29), .Cin(c_28_28));
    full_adder adder_28_30(.S(s_28_30), .Cout(c_28_30), .A(s_27_30), .B(w_28_30), .Cin(c_28_29));
    full_adder adder_28_31(.S(s_28_31), .Cout(c_28_31), .A(s_27_31), .B(w_28_31), .Cin(c_28_30));
    full_adder adder_28_32(.S(s_28_32), .Cout(c_28_32), .A(s_27_32), .B(w_28_32), .Cin(c_28_31));
    full_adder adder_28_33(.S(s_28_33), .Cout(c_28_33), .A(s_27_33), .B(w_28_33), .Cin(c_28_32));
    full_adder adder_28_34(.S(s_28_34), .Cout(c_28_34), .A(s_27_34), .B(w_28_34), .Cin(c_28_33));
    full_adder adder_28_35(.S(s_28_35), .Cout(c_28_35), .A(s_27_35), .B(w_28_35), .Cin(c_28_34));
    full_adder adder_28_36(.S(s_28_36), .Cout(c_28_36), .A(s_27_36), .B(w_28_36), .Cin(c_28_35));
    full_adder adder_28_37(.S(s_28_37), .Cout(c_28_37), .A(s_27_37), .B(w_28_37), .Cin(c_28_36));
    full_adder adder_28_38(.S(s_28_38), .Cout(c_28_38), .A(s_27_38), .B(w_28_38), .Cin(c_28_37));
    full_adder adder_28_39(.S(s_28_39), .Cout(c_28_39), .A(s_27_39), .B(w_28_39), .Cin(c_28_38));
    full_adder adder_28_40(.S(s_28_40), .Cout(c_28_40), .A(s_27_40), .B(w_28_40), .Cin(c_28_39));
    full_adder adder_28_41(.S(s_28_41), .Cout(c_28_41), .A(s_27_41), .B(w_28_41), .Cin(c_28_40));
    full_adder adder_28_42(.S(s_28_42), .Cout(c_28_42), .A(s_27_42), .B(w_28_42), .Cin(c_28_41));
    full_adder adder_28_43(.S(s_28_43), .Cout(c_28_43), .A(s_27_43), .B(w_28_43), .Cin(c_28_42));
    full_adder adder_28_44(.S(s_28_44), .Cout(c_28_44), .A(s_27_44), .B(w_28_44), .Cin(c_28_43));
    full_adder adder_28_45(.S(s_28_45), .Cout(c_28_45), .A(s_27_45), .B(w_28_45), .Cin(c_28_44));
    full_adder adder_28_46(.S(s_28_46), .Cout(c_28_46), .A(s_27_46), .B(w_28_46), .Cin(c_28_45));
    full_adder adder_28_47(.S(s_28_47), .Cout(c_28_47), .A(s_27_47), .B(w_28_47), .Cin(c_28_46));
    full_adder adder_28_48(.S(s_28_48), .Cout(c_28_48), .A(s_27_48), .B(w_28_48), .Cin(c_28_47));
    full_adder adder_28_49(.S(s_28_49), .Cout(c_28_49), .A(s_27_49), .B(w_28_49), .Cin(c_28_48));
    full_adder adder_28_50(.S(s_28_50), .Cout(c_28_50), .A(s_27_50), .B(w_28_50), .Cin(c_28_49));
    full_adder adder_28_51(.S(s_28_51), .Cout(c_28_51), .A(s_27_51), .B(w_28_51), .Cin(c_28_50));
    full_adder adder_28_52(.S(s_28_52), .Cout(c_28_52), .A(s_27_52), .B(w_28_52), .Cin(c_28_51));
    full_adder adder_28_53(.S(s_28_53), .Cout(c_28_53), .A(s_27_53), .B(w_28_53), .Cin(c_28_52));
    full_adder adder_28_54(.S(s_28_54), .Cout(c_28_54), .A(s_27_54), .B(w_28_54), .Cin(c_28_53));
    full_adder adder_28_55(.S(s_28_55), .Cout(c_28_55), .A(s_27_55), .B(w_28_55), .Cin(c_28_54));
    full_adder adder_28_56(.S(s_28_56), .Cout(c_28_56), .A(s_27_56), .B(w_28_56), .Cin(c_28_55));
    full_adder adder_28_57(.S(s_28_57), .Cout(c_28_57), .A(s_27_57), .B(w_28_57), .Cin(c_28_56));
    full_adder adder_28_58(.S(s_28_58), .Cout(c_28_58), .A(s_27_58), .B(w_28_58), .Cin(c_28_57));
    full_adder adder_28_59(.S(s_28_59), .Cout(c_28_59), .A(c_27_58), .B(w_28_59), .Cin(c_28_58));
    assign result[28] = s_28_28;
    wire w_29_29, w_29_30, w_29_31, w_29_32, w_29_33, w_29_34, w_29_35, w_29_36, w_29_37, w_29_38, w_29_39, w_29_40, w_29_41, w_29_42, w_29_43, w_29_44, w_29_45, w_29_46, w_29_47, w_29_48, w_29_49, w_29_50, w_29_51, w_29_52, w_29_53, w_29_54, w_29_55, w_29_56, w_29_57, w_29_58, w_29_59, w_29_60;
    wire s_29_29, s_29_30, s_29_31, s_29_32, s_29_33, s_29_34, s_29_35, s_29_36, s_29_37, s_29_38, s_29_39, s_29_40, s_29_41, s_29_42, s_29_43, s_29_44, s_29_45, s_29_46, s_29_47, s_29_48, s_29_49, s_29_50, s_29_51, s_29_52, s_29_53, s_29_54, s_29_55, s_29_56, s_29_57, s_29_58, s_29_59, s_29_60;
    wire c_29_29, c_29_30, c_29_31, c_29_32, c_29_33, c_29_34, c_29_35, c_29_36, c_29_37, c_29_38, c_29_39, c_29_40, c_29_41, c_29_42, c_29_43, c_29_44, c_29_45, c_29_46, c_29_47, c_29_48, c_29_49, c_29_50, c_29_51, c_29_52, c_29_53, c_29_54, c_29_55, c_29_56, c_29_57, c_29_58, c_29_59, c_29_60;
    assign w_29_29 = data_operandA[0] & data_operandB[29];
    assign w_29_30 = data_operandA[1] & data_operandB[29];
    assign w_29_31 = data_operandA[2] & data_operandB[29];
    assign w_29_32 = data_operandA[3] & data_operandB[29];
    assign w_29_33 = data_operandA[4] & data_operandB[29];
    assign w_29_34 = data_operandA[5] & data_operandB[29];
    assign w_29_35 = data_operandA[6] & data_operandB[29];
    assign w_29_36 = data_operandA[7] & data_operandB[29];
    assign w_29_37 = data_operandA[8] & data_operandB[29];
    assign w_29_38 = data_operandA[9] & data_operandB[29];
    assign w_29_39 = data_operandA[10] & data_operandB[29];
    assign w_29_40 = data_operandA[11] & data_operandB[29];
    assign w_29_41 = data_operandA[12] & data_operandB[29];
    assign w_29_42 = data_operandA[13] & data_operandB[29];
    assign w_29_43 = data_operandA[14] & data_operandB[29];
    assign w_29_44 = data_operandA[15] & data_operandB[29];
    assign w_29_45 = data_operandA[16] & data_operandB[29];
    assign w_29_46 = data_operandA[17] & data_operandB[29];
    assign w_29_47 = data_operandA[18] & data_operandB[29];
    assign w_29_48 = data_operandA[19] & data_operandB[29];
    assign w_29_49 = data_operandA[20] & data_operandB[29];
    assign w_29_50 = data_operandA[21] & data_operandB[29];
    assign w_29_51 = data_operandA[22] & data_operandB[29];
    assign w_29_52 = data_operandA[23] & data_operandB[29];
    assign w_29_53 = data_operandA[24] & data_operandB[29];
    assign w_29_54 = data_operandA[25] & data_operandB[29];
    assign w_29_55 = data_operandA[26] & data_operandB[29];
    assign w_29_56 = data_operandA[27] & data_operandB[29];
    assign w_29_57 = data_operandA[28] & data_operandB[29];
    assign w_29_58 = data_operandA[29] & data_operandB[29];
    assign w_29_59 = data_operandA[30] & data_operandB[29];
    assign w_29_60 = ~(data_operandA[31] & data_operandB[29]);
    full_adder adder_29_29(.S(s_29_29), .Cout(c_29_29), .A(s_28_29), .B(w_29_29), .Cin(1'b0));
    full_adder adder_29_30(.S(s_29_30), .Cout(c_29_30), .A(s_28_30), .B(w_29_30), .Cin(c_29_29));
    full_adder adder_29_31(.S(s_29_31), .Cout(c_29_31), .A(s_28_31), .B(w_29_31), .Cin(c_29_30));
    full_adder adder_29_32(.S(s_29_32), .Cout(c_29_32), .A(s_28_32), .B(w_29_32), .Cin(c_29_31));
    full_adder adder_29_33(.S(s_29_33), .Cout(c_29_33), .A(s_28_33), .B(w_29_33), .Cin(c_29_32));
    full_adder adder_29_34(.S(s_29_34), .Cout(c_29_34), .A(s_28_34), .B(w_29_34), .Cin(c_29_33));
    full_adder adder_29_35(.S(s_29_35), .Cout(c_29_35), .A(s_28_35), .B(w_29_35), .Cin(c_29_34));
    full_adder adder_29_36(.S(s_29_36), .Cout(c_29_36), .A(s_28_36), .B(w_29_36), .Cin(c_29_35));
    full_adder adder_29_37(.S(s_29_37), .Cout(c_29_37), .A(s_28_37), .B(w_29_37), .Cin(c_29_36));
    full_adder adder_29_38(.S(s_29_38), .Cout(c_29_38), .A(s_28_38), .B(w_29_38), .Cin(c_29_37));
    full_adder adder_29_39(.S(s_29_39), .Cout(c_29_39), .A(s_28_39), .B(w_29_39), .Cin(c_29_38));
    full_adder adder_29_40(.S(s_29_40), .Cout(c_29_40), .A(s_28_40), .B(w_29_40), .Cin(c_29_39));
    full_adder adder_29_41(.S(s_29_41), .Cout(c_29_41), .A(s_28_41), .B(w_29_41), .Cin(c_29_40));
    full_adder adder_29_42(.S(s_29_42), .Cout(c_29_42), .A(s_28_42), .B(w_29_42), .Cin(c_29_41));
    full_adder adder_29_43(.S(s_29_43), .Cout(c_29_43), .A(s_28_43), .B(w_29_43), .Cin(c_29_42));
    full_adder adder_29_44(.S(s_29_44), .Cout(c_29_44), .A(s_28_44), .B(w_29_44), .Cin(c_29_43));
    full_adder adder_29_45(.S(s_29_45), .Cout(c_29_45), .A(s_28_45), .B(w_29_45), .Cin(c_29_44));
    full_adder adder_29_46(.S(s_29_46), .Cout(c_29_46), .A(s_28_46), .B(w_29_46), .Cin(c_29_45));
    full_adder adder_29_47(.S(s_29_47), .Cout(c_29_47), .A(s_28_47), .B(w_29_47), .Cin(c_29_46));
    full_adder adder_29_48(.S(s_29_48), .Cout(c_29_48), .A(s_28_48), .B(w_29_48), .Cin(c_29_47));
    full_adder adder_29_49(.S(s_29_49), .Cout(c_29_49), .A(s_28_49), .B(w_29_49), .Cin(c_29_48));
    full_adder adder_29_50(.S(s_29_50), .Cout(c_29_50), .A(s_28_50), .B(w_29_50), .Cin(c_29_49));
    full_adder adder_29_51(.S(s_29_51), .Cout(c_29_51), .A(s_28_51), .B(w_29_51), .Cin(c_29_50));
    full_adder adder_29_52(.S(s_29_52), .Cout(c_29_52), .A(s_28_52), .B(w_29_52), .Cin(c_29_51));
    full_adder adder_29_53(.S(s_29_53), .Cout(c_29_53), .A(s_28_53), .B(w_29_53), .Cin(c_29_52));
    full_adder adder_29_54(.S(s_29_54), .Cout(c_29_54), .A(s_28_54), .B(w_29_54), .Cin(c_29_53));
    full_adder adder_29_55(.S(s_29_55), .Cout(c_29_55), .A(s_28_55), .B(w_29_55), .Cin(c_29_54));
    full_adder adder_29_56(.S(s_29_56), .Cout(c_29_56), .A(s_28_56), .B(w_29_56), .Cin(c_29_55));
    full_adder adder_29_57(.S(s_29_57), .Cout(c_29_57), .A(s_28_57), .B(w_29_57), .Cin(c_29_56));
    full_adder adder_29_58(.S(s_29_58), .Cout(c_29_58), .A(s_28_58), .B(w_29_58), .Cin(c_29_57));
    full_adder adder_29_59(.S(s_29_59), .Cout(c_29_59), .A(s_28_59), .B(w_29_59), .Cin(c_29_58));
    full_adder adder_29_60(.S(s_29_60), .Cout(c_29_60), .A(c_28_59), .B(w_29_60), .Cin(c_29_59));
    assign result[29] = s_29_29;
    wire w_30_30, w_30_31, w_30_32, w_30_33, w_30_34, w_30_35, w_30_36, w_30_37, w_30_38, w_30_39, w_30_40, w_30_41, w_30_42, w_30_43, w_30_44, w_30_45, w_30_46, w_30_47, w_30_48, w_30_49, w_30_50, w_30_51, w_30_52, w_30_53, w_30_54, w_30_55, w_30_56, w_30_57, w_30_58, w_30_59, w_30_60, w_30_61;
    wire s_30_30, s_30_31, s_30_32, s_30_33, s_30_34, s_30_35, s_30_36, s_30_37, s_30_38, s_30_39, s_30_40, s_30_41, s_30_42, s_30_43, s_30_44, s_30_45, s_30_46, s_30_47, s_30_48, s_30_49, s_30_50, s_30_51, s_30_52, s_30_53, s_30_54, s_30_55, s_30_56, s_30_57, s_30_58, s_30_59, s_30_60, s_30_61;
    wire c_30_30, c_30_31, c_30_32, c_30_33, c_30_34, c_30_35, c_30_36, c_30_37, c_30_38, c_30_39, c_30_40, c_30_41, c_30_42, c_30_43, c_30_44, c_30_45, c_30_46, c_30_47, c_30_48, c_30_49, c_30_50, c_30_51, c_30_52, c_30_53, c_30_54, c_30_55, c_30_56, c_30_57, c_30_58, c_30_59, c_30_60, c_30_61;
    assign w_30_30 = data_operandA[0] & data_operandB[30];
    assign w_30_31 = data_operandA[1] & data_operandB[30];
    assign w_30_32 = data_operandA[2] & data_operandB[30];
    assign w_30_33 = data_operandA[3] & data_operandB[30];
    assign w_30_34 = data_operandA[4] & data_operandB[30];
    assign w_30_35 = data_operandA[5] & data_operandB[30];
    assign w_30_36 = data_operandA[6] & data_operandB[30];
    assign w_30_37 = data_operandA[7] & data_operandB[30];
    assign w_30_38 = data_operandA[8] & data_operandB[30];
    assign w_30_39 = data_operandA[9] & data_operandB[30];
    assign w_30_40 = data_operandA[10] & data_operandB[30];
    assign w_30_41 = data_operandA[11] & data_operandB[30];
    assign w_30_42 = data_operandA[12] & data_operandB[30];
    assign w_30_43 = data_operandA[13] & data_operandB[30];
    assign w_30_44 = data_operandA[14] & data_operandB[30];
    assign w_30_45 = data_operandA[15] & data_operandB[30];
    assign w_30_46 = data_operandA[16] & data_operandB[30];
    assign w_30_47 = data_operandA[17] & data_operandB[30];
    assign w_30_48 = data_operandA[18] & data_operandB[30];
    assign w_30_49 = data_operandA[19] & data_operandB[30];
    assign w_30_50 = data_operandA[20] & data_operandB[30];
    assign w_30_51 = data_operandA[21] & data_operandB[30];
    assign w_30_52 = data_operandA[22] & data_operandB[30];
    assign w_30_53 = data_operandA[23] & data_operandB[30];
    assign w_30_54 = data_operandA[24] & data_operandB[30];
    assign w_30_55 = data_operandA[25] & data_operandB[30];
    assign w_30_56 = data_operandA[26] & data_operandB[30];
    assign w_30_57 = data_operandA[27] & data_operandB[30];
    assign w_30_58 = data_operandA[28] & data_operandB[30];
    assign w_30_59 = data_operandA[29] & data_operandB[30];
    assign w_30_60 = data_operandA[30] & data_operandB[30];
    assign w_30_61 = ~(data_operandA[31] & data_operandB[30]);
    full_adder adder_30_30(.S(s_30_30), .Cout(c_30_30), .A(s_29_30), .B(w_30_30), .Cin(1'b0));
    full_adder adder_30_31(.S(s_30_31), .Cout(c_30_31), .A(s_29_31), .B(w_30_31), .Cin(c_30_30));
    full_adder adder_30_32(.S(s_30_32), .Cout(c_30_32), .A(s_29_32), .B(w_30_32), .Cin(c_30_31));
    full_adder adder_30_33(.S(s_30_33), .Cout(c_30_33), .A(s_29_33), .B(w_30_33), .Cin(c_30_32));
    full_adder adder_30_34(.S(s_30_34), .Cout(c_30_34), .A(s_29_34), .B(w_30_34), .Cin(c_30_33));
    full_adder adder_30_35(.S(s_30_35), .Cout(c_30_35), .A(s_29_35), .B(w_30_35), .Cin(c_30_34));
    full_adder adder_30_36(.S(s_30_36), .Cout(c_30_36), .A(s_29_36), .B(w_30_36), .Cin(c_30_35));
    full_adder adder_30_37(.S(s_30_37), .Cout(c_30_37), .A(s_29_37), .B(w_30_37), .Cin(c_30_36));
    full_adder adder_30_38(.S(s_30_38), .Cout(c_30_38), .A(s_29_38), .B(w_30_38), .Cin(c_30_37));
    full_adder adder_30_39(.S(s_30_39), .Cout(c_30_39), .A(s_29_39), .B(w_30_39), .Cin(c_30_38));
    full_adder adder_30_40(.S(s_30_40), .Cout(c_30_40), .A(s_29_40), .B(w_30_40), .Cin(c_30_39));
    full_adder adder_30_41(.S(s_30_41), .Cout(c_30_41), .A(s_29_41), .B(w_30_41), .Cin(c_30_40));
    full_adder adder_30_42(.S(s_30_42), .Cout(c_30_42), .A(s_29_42), .B(w_30_42), .Cin(c_30_41));
    full_adder adder_30_43(.S(s_30_43), .Cout(c_30_43), .A(s_29_43), .B(w_30_43), .Cin(c_30_42));
    full_adder adder_30_44(.S(s_30_44), .Cout(c_30_44), .A(s_29_44), .B(w_30_44), .Cin(c_30_43));
    full_adder adder_30_45(.S(s_30_45), .Cout(c_30_45), .A(s_29_45), .B(w_30_45), .Cin(c_30_44));
    full_adder adder_30_46(.S(s_30_46), .Cout(c_30_46), .A(s_29_46), .B(w_30_46), .Cin(c_30_45));
    full_adder adder_30_47(.S(s_30_47), .Cout(c_30_47), .A(s_29_47), .B(w_30_47), .Cin(c_30_46));
    full_adder adder_30_48(.S(s_30_48), .Cout(c_30_48), .A(s_29_48), .B(w_30_48), .Cin(c_30_47));
    full_adder adder_30_49(.S(s_30_49), .Cout(c_30_49), .A(s_29_49), .B(w_30_49), .Cin(c_30_48));
    full_adder adder_30_50(.S(s_30_50), .Cout(c_30_50), .A(s_29_50), .B(w_30_50), .Cin(c_30_49));
    full_adder adder_30_51(.S(s_30_51), .Cout(c_30_51), .A(s_29_51), .B(w_30_51), .Cin(c_30_50));
    full_adder adder_30_52(.S(s_30_52), .Cout(c_30_52), .A(s_29_52), .B(w_30_52), .Cin(c_30_51));
    full_adder adder_30_53(.S(s_30_53), .Cout(c_30_53), .A(s_29_53), .B(w_30_53), .Cin(c_30_52));
    full_adder adder_30_54(.S(s_30_54), .Cout(c_30_54), .A(s_29_54), .B(w_30_54), .Cin(c_30_53));
    full_adder adder_30_55(.S(s_30_55), .Cout(c_30_55), .A(s_29_55), .B(w_30_55), .Cin(c_30_54));
    full_adder adder_30_56(.S(s_30_56), .Cout(c_30_56), .A(s_29_56), .B(w_30_56), .Cin(c_30_55));
    full_adder adder_30_57(.S(s_30_57), .Cout(c_30_57), .A(s_29_57), .B(w_30_57), .Cin(c_30_56));
    full_adder adder_30_58(.S(s_30_58), .Cout(c_30_58), .A(s_29_58), .B(w_30_58), .Cin(c_30_57));
    full_adder adder_30_59(.S(s_30_59), .Cout(c_30_59), .A(s_29_59), .B(w_30_59), .Cin(c_30_58));
    full_adder adder_30_60(.S(s_30_60), .Cout(c_30_60), .A(s_29_60), .B(w_30_60), .Cin(c_30_59));
    full_adder adder_30_61(.S(s_30_61), .Cout(c_30_61), .A(c_29_60), .B(w_30_61), .Cin(c_30_60));
    assign result[30] = s_30_30;
    wire w_31_31, w_31_32, w_31_33, w_31_34, w_31_35, w_31_36, w_31_37, w_31_38, w_31_39, w_31_40, w_31_41, w_31_42, w_31_43, w_31_44, w_31_45, w_31_46, w_31_47, w_31_48, w_31_49, w_31_50, w_31_51, w_31_52, w_31_53, w_31_54, w_31_55, w_31_56, w_31_57, w_31_58, w_31_59, w_31_60, w_31_61, w_31_62;
    wire s_31_31, s_31_32, s_31_33, s_31_34, s_31_35, s_31_36, s_31_37, s_31_38, s_31_39, s_31_40, s_31_41, s_31_42, s_31_43, s_31_44, s_31_45, s_31_46, s_31_47, s_31_48, s_31_49, s_31_50, s_31_51, s_31_52, s_31_53, s_31_54, s_31_55, s_31_56, s_31_57, s_31_58, s_31_59, s_31_60, s_31_61, s_31_62;
    wire s_31_63;
    wire c_31_31, c_31_32, c_31_33, c_31_34, c_31_35, c_31_36, c_31_37, c_31_38, c_31_39, c_31_40, c_31_41, c_31_42, c_31_43, c_31_44, c_31_45, c_31_46, c_31_47, c_31_48, c_31_49, c_31_50, c_31_51, c_31_52, c_31_53, c_31_54, c_31_55, c_31_56, c_31_57, c_31_58, c_31_59, c_31_60, c_31_61, c_31_62;
    wire c_31_63;
    assign w_31_31 = ~(data_operandA[0] & data_operandB[31]);
    assign w_31_32 = ~(data_operandA[1] & data_operandB[31]);
    assign w_31_33 = ~(data_operandA[2] & data_operandB[31]);
    assign w_31_34 = ~(data_operandA[3] & data_operandB[31]);
    assign w_31_35 = ~(data_operandA[4] & data_operandB[31]);
    assign w_31_36 = ~(data_operandA[5] & data_operandB[31]);
    assign w_31_37 = ~(data_operandA[6] & data_operandB[31]);
    assign w_31_38 = ~(data_operandA[7] & data_operandB[31]);
    assign w_31_39 = ~(data_operandA[8] & data_operandB[31]);
    assign w_31_40 = ~(data_operandA[9] & data_operandB[31]);
    assign w_31_41 = ~(data_operandA[10] & data_operandB[31]);
    assign w_31_42 = ~(data_operandA[11] & data_operandB[31]);
    assign w_31_43 = ~(data_operandA[12] & data_operandB[31]);
    assign w_31_44 = ~(data_operandA[13] & data_operandB[31]);
    assign w_31_45 = ~(data_operandA[14] & data_operandB[31]);
    assign w_31_46 = ~(data_operandA[15] & data_operandB[31]);
    assign w_31_47 = ~(data_operandA[16] & data_operandB[31]);
    assign w_31_48 = ~(data_operandA[17] & data_operandB[31]);
    assign w_31_49 = ~(data_operandA[18] & data_operandB[31]);
    assign w_31_50 = ~(data_operandA[19] & data_operandB[31]);
    assign w_31_51 = ~(data_operandA[20] & data_operandB[31]);
    assign w_31_52 = ~(data_operandA[21] & data_operandB[31]);
    assign w_31_53 = ~(data_operandA[22] & data_operandB[31]);
    assign w_31_54 = ~(data_operandA[23] & data_operandB[31]);
    assign w_31_55 = ~(data_operandA[24] & data_operandB[31]);
    assign w_31_56 = ~(data_operandA[25] & data_operandB[31]);
    assign w_31_57 = ~(data_operandA[26] & data_operandB[31]);
    assign w_31_58 = ~(data_operandA[27] & data_operandB[31]);
    assign w_31_59 = ~(data_operandA[28] & data_operandB[31]);
    assign w_31_60 = ~(data_operandA[29] & data_operandB[31]);
    assign w_31_61 = ~(data_operandA[30] & data_operandB[31]);
    assign w_31_62 = data_operandA[31] & data_operandB[31];
    full_adder adder_31_31(.S(s_31_31), .Cout(c_31_31), .A(s_30_31), .B(w_31_31), .Cin(1'b0));
    full_adder adder_31_32(.S(s_31_32), .Cout(c_31_32), .A(s_30_32), .B(w_31_32), .Cin(c_31_31));
    full_adder adder_31_33(.S(s_31_33), .Cout(c_31_33), .A(s_30_33), .B(w_31_33), .Cin(c_31_32));
    full_adder adder_31_34(.S(s_31_34), .Cout(c_31_34), .A(s_30_34), .B(w_31_34), .Cin(c_31_33));
    full_adder adder_31_35(.S(s_31_35), .Cout(c_31_35), .A(s_30_35), .B(w_31_35), .Cin(c_31_34));
    full_adder adder_31_36(.S(s_31_36), .Cout(c_31_36), .A(s_30_36), .B(w_31_36), .Cin(c_31_35));
    full_adder adder_31_37(.S(s_31_37), .Cout(c_31_37), .A(s_30_37), .B(w_31_37), .Cin(c_31_36));
    full_adder adder_31_38(.S(s_31_38), .Cout(c_31_38), .A(s_30_38), .B(w_31_38), .Cin(c_31_37));
    full_adder adder_31_39(.S(s_31_39), .Cout(c_31_39), .A(s_30_39), .B(w_31_39), .Cin(c_31_38));
    full_adder adder_31_40(.S(s_31_40), .Cout(c_31_40), .A(s_30_40), .B(w_31_40), .Cin(c_31_39));
    full_adder adder_31_41(.S(s_31_41), .Cout(c_31_41), .A(s_30_41), .B(w_31_41), .Cin(c_31_40));
    full_adder adder_31_42(.S(s_31_42), .Cout(c_31_42), .A(s_30_42), .B(w_31_42), .Cin(c_31_41));
    full_adder adder_31_43(.S(s_31_43), .Cout(c_31_43), .A(s_30_43), .B(w_31_43), .Cin(c_31_42));
    full_adder adder_31_44(.S(s_31_44), .Cout(c_31_44), .A(s_30_44), .B(w_31_44), .Cin(c_31_43));
    full_adder adder_31_45(.S(s_31_45), .Cout(c_31_45), .A(s_30_45), .B(w_31_45), .Cin(c_31_44));
    full_adder adder_31_46(.S(s_31_46), .Cout(c_31_46), .A(s_30_46), .B(w_31_46), .Cin(c_31_45));
    full_adder adder_31_47(.S(s_31_47), .Cout(c_31_47), .A(s_30_47), .B(w_31_47), .Cin(c_31_46));
    full_adder adder_31_48(.S(s_31_48), .Cout(c_31_48), .A(s_30_48), .B(w_31_48), .Cin(c_31_47));
    full_adder adder_31_49(.S(s_31_49), .Cout(c_31_49), .A(s_30_49), .B(w_31_49), .Cin(c_31_48));
    full_adder adder_31_50(.S(s_31_50), .Cout(c_31_50), .A(s_30_50), .B(w_31_50), .Cin(c_31_49));
    full_adder adder_31_51(.S(s_31_51), .Cout(c_31_51), .A(s_30_51), .B(w_31_51), .Cin(c_31_50));
    full_adder adder_31_52(.S(s_31_52), .Cout(c_31_52), .A(s_30_52), .B(w_31_52), .Cin(c_31_51));
    full_adder adder_31_53(.S(s_31_53), .Cout(c_31_53), .A(s_30_53), .B(w_31_53), .Cin(c_31_52));
    full_adder adder_31_54(.S(s_31_54), .Cout(c_31_54), .A(s_30_54), .B(w_31_54), .Cin(c_31_53));
    full_adder adder_31_55(.S(s_31_55), .Cout(c_31_55), .A(s_30_55), .B(w_31_55), .Cin(c_31_54));
    full_adder adder_31_56(.S(s_31_56), .Cout(c_31_56), .A(s_30_56), .B(w_31_56), .Cin(c_31_55));
    full_adder adder_31_57(.S(s_31_57), .Cout(c_31_57), .A(s_30_57), .B(w_31_57), .Cin(c_31_56));
    full_adder adder_31_58(.S(s_31_58), .Cout(c_31_58), .A(s_30_58), .B(w_31_58), .Cin(c_31_57));
    full_adder adder_31_59(.S(s_31_59), .Cout(c_31_59), .A(s_30_59), .B(w_31_59), .Cin(c_31_58));
    full_adder adder_31_60(.S(s_31_60), .Cout(c_31_60), .A(s_30_60), .B(w_31_60), .Cin(c_31_59));
    full_adder adder_31_61(.S(s_31_61), .Cout(c_31_61), .A(s_30_61), .B(w_31_61), .Cin(c_31_60));
    full_adder adder_31_62(.S(s_31_62), .Cout(c_31_62), .A(c_30_61), .B(w_31_62), .Cin(c_31_61));
    full_adder adder_31_63(.S(s_31_63), .Cout(c_31_63), .A(1'b1), .B(c_31_62), .Cin(1'b0));
    assign result[31] = s_31_31;
    assign result[32] = s_31_32;
    assign result[33] = s_31_33;
    assign result[34] = s_31_34;
    assign result[35] = s_31_35;
    assign result[36] = s_31_36;
    assign result[37] = s_31_37;
    assign result[38] = s_31_38;
    assign result[39] = s_31_39;
    assign result[40] = s_31_40;
    assign result[41] = s_31_41;
    assign result[42] = s_31_42;
    assign result[43] = s_31_43;
    assign result[44] = s_31_44;
    assign result[45] = s_31_45;
    assign result[46] = s_31_46;
    assign result[47] = s_31_47;
    assign result[48] = s_31_48;
    assign result[49] = s_31_49;
    assign result[50] = s_31_50;
    assign result[51] = s_31_51;
    assign result[52] = s_31_52;
    assign result[53] = s_31_53;
    assign result[54] = s_31_54;
    assign result[55] = s_31_55;
    assign result[56] = s_31_56;
    assign result[57] = s_31_57;
    assign result[58] = s_31_58;
    assign result[59] = s_31_59;
    assign result[60] = s_31_60;
    assign result[61] = s_31_61;
    assign result[62] = s_31_62;
    assign result[63] = s_31_63;

endmodule