module sr_4b(out, data_operandA);

    input [31:0] data_operandA;
    output [31:0] out;

    assign out[0] = data_operandA[4];
    assign out[1] = data_operandA[5];
    assign out[2] = data_operandA[6];
    assign out[3] = data_operandA[7];
    assign out[4] = data_operandA[8];
    assign out[5] = data_operandA[9];
    assign out[6] = data_operandA[10];
    assign out[7] = data_operandA[11];
    assign out[8] = data_operandA[12];
    assign out[9] = data_operandA[13];
    assign out[10] = data_operandA[14];
    assign out[11] = data_operandA[15];
    assign out[12] = data_operandA[16];
    assign out[13] = data_operandA[17];
    assign out[14] = data_operandA[18];
    assign out[15] = data_operandA[19];
    assign out[16] = data_operandA[20];
    assign out[17] = data_operandA[21];
    assign out[18] = data_operandA[22];
    assign out[19] = data_operandA[23];
    assign out[20] = data_operandA[24];
    assign out[21] = data_operandA[25];
    assign out[22] = data_operandA[26];
    assign out[23] = data_operandA[27];
    assign out[24] = data_operandA[28];
    assign out[25] = data_operandA[29];
    assign out[26] = data_operandA[30];
    assign out[27] = data_operandA[31];
    assign out[28] = data_operandA[31];
    assign out[29] = data_operandA[31];
    assign out[30] = data_operandA[31];
    assign out[31] = data_operandA[31];


endmodule