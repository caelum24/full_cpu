module and_32bit(result, A, B);

    input [31:0] A, B;
    output [31:0] result;

    and a0(result[0], A[0], B[0]);
    and a1(result[1], A[1], B[1]);
    and a2(result[2], A[2], B[2]);
    and a3(result[3], A[3], B[3]);
    and a4(result[4], A[4], B[4]);
    and a5(result[5], A[5], B[5]);
    and a6(result[6], A[6], B[6]);
    and a7(result[7], A[7], B[7]);
    and a8(result[8], A[8], B[8]);
    and a9(result[9], A[9], B[9]);
    and a10(result[10], A[10], B[10]);
    and a11(result[11], A[11], B[11]);
    and a12(result[12], A[12], B[12]);
    and a13(result[13], A[13], B[13]);
    and a14(result[14], A[14], B[14]);
    and a15(result[15], A[15], B[15]);
    and a16(result[16], A[16], B[16]);
    and a17(result[17], A[17], B[17]);
    and a18(result[18], A[18], B[18]);
    and a19(result[19], A[19], B[19]);
    and a20(result[20], A[20], B[20]);
    and a21(result[21], A[21], B[21]);
    and a22(result[22], A[22], B[22]);
    and a23(result[23], A[23], B[23]);
    and a24(result[24], A[24], B[24]);
    and a25(result[25], A[25], B[25]);
    and a26(result[26], A[26], B[26]);
    and a27(result[27], A[27], B[27]);
    and a28(result[28], A[28], B[28]);
    and a29(result[29], A[29], B[29]);
    and a30(result[30], A[30], B[30]);
    and a31(result[31], A[31], B[31]);

endmodule